module HRALM4 (clk,
    rst,
    p,
    x,
    y);
 input clk;
 input rst;
 output [31:0] p;
 input [15:0] x;
 input [15:0] y;

 wire \ADDER.A1.Sum[0] ;
 wire \ADDER.A4.Sum[0] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire net62;
 wire _0117_;
 wire net61;
 wire net60;
 wire net59;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire net58;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire net57;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire net55;
 wire net54;
 wire _0137_;
 wire net53;
 wire net52;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire net51;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire net50;
 wire _0152_;
 wire _0153_;
 wire net49;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire net48;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire net46;
 wire _0189_;
 wire net45;
 wire net44;
 wire _0192_;
 wire _0193_;
 wire net43;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire net42;
 wire net41;
 wire _0217_;
 wire net40;
 wire net39;
 wire net38;
 wire _0221_;
 wire net37;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire net36;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire net35;
 wire _0235_;
 wire net34;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire net33;
 wire _0243_;
 wire net32;
 wire _0245_;
 wire net31;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire net30;
 wire net29;
 wire net28;
 wire _0255_;
 wire net27;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire net26;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire net25;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire net24;
 wire net23;
 wire _0287_;
 wire _0288_;
 wire net22;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire net21;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire net20;
 wire net19;
 wire net18;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire net17;
 wire _0363_;
 wire _0364_;
 wire net16;
 wire _0366_;
 wire net15;
 wire net14;
 wire net13;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire net12;
 wire _0382_;
 wire net11;
 wire net10;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire net9;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire net8;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire net6;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire net5;
 wire _0529_;
 wire net4;
 wire net3;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire net2;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire net1;
 wire _0621_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire net47;
 wire _0692_;
 wire _0693_;
 wire net56;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire net7;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire \add1.sm ;
 wire net63;
 wire net64;
 wire net65;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;

 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_63 ();
 INVx1_ASAP7_75t_R _0754_ (.A(net3),
    .Y(_0117_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_60 ();
 OR2x2_ASAP7_75t_R _0758_ (.A(net5),
    .B(net172),
    .Y(_0121_));
 OR3x1_ASAP7_75t_R _0759_ (.A(_0117_),
    .B(net4),
    .C(_0121_),
    .Y(_0122_));
 INVx3_ASAP7_75t_R _0760_ (.A(net4),
    .Y(_0123_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_59 ();
 NAND2x2_ASAP7_75t_R _0762_ (.A(net5),
    .B(net176),
    .Y(_0125_));
 OR3x1_ASAP7_75t_R _0763_ (.A(net3),
    .B(_0123_),
    .C(_0125_),
    .Y(_0126_));
 INVx1_ASAP7_75t_R _0764_ (.A(net16),
    .Y(_0127_));
 NOR2x1_ASAP7_75t_R _0765_ (.A(net5),
    .B(net176),
    .Y(_0128_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_58 ();
 NOR3x1_ASAP7_75t_R _0767_ (.A(net17),
    .B(net3),
    .C(net4),
    .Y(_0130_));
 AND4x1_ASAP7_75t_R _0768_ (.A(net16),
    .B(net17),
    .C(net3),
    .D(net4),
    .Y(_0131_));
 AND2x2_ASAP7_75t_R _0769_ (.A(net6),
    .B(net5),
    .Y(_0132_));
 AO32x2_ASAP7_75t_R _0770_ (.A1(_0127_),
    .A2(_0128_),
    .A3(_0130_),
    .B1(_0131_),
    .B2(_0132_),
    .Y(_0133_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_57 ();
 INVx2_ASAP7_75t_R _0772_ (.A(net95),
    .Y(_0134_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_55 ();
 NAND3x2_ASAP7_75t_R _0775_ (.B(net14),
    .C(net15),
    .Y(_0137_),
    .A(net6));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_53 ();
 NAND2x1_ASAP7_75t_R _0778_ (.A(net12),
    .B(net13),
    .Y(_0140_));
 OR5x1_ASAP7_75t_R _0779_ (.A(net6),
    .B(net12),
    .C(net13),
    .D(net14),
    .E(net15),
    .Y(_0141_));
 OA21x2_ASAP7_75t_R _0780_ (.A1(_0137_),
    .A2(_0140_),
    .B(_0141_),
    .Y(_0142_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_52 ();
 INVx2_ASAP7_75t_R _0782_ (.A(net11),
    .Y(_0144_));
 NAND2x1_ASAP7_75t_R _0783_ (.A(net10),
    .B(_0144_),
    .Y(_0145_));
 CKINVDCx5p33_ASAP7_75t_R _0784_ (.A(net176),
    .Y(_0146_));
 INVx5_ASAP7_75t_R _0785_ (.A(net15),
    .Y(_0147_));
 NAND2x1_ASAP7_75t_R _0786_ (.A(net14),
    .B(_0147_),
    .Y(_0148_));
 OA211x2_ASAP7_75t_R _0787_ (.A1(_0142_),
    .A2(_0145_),
    .B(_0146_),
    .C(_0148_),
    .Y(_0149_));
 INVx2_ASAP7_75t_R _0788_ (.A(net10),
    .Y(_0150_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Right_51 ();
 NAND2x1_ASAP7_75t_R _0790_ (.A(_0150_),
    .B(net11),
    .Y(_0152_));
 INVx2_ASAP7_75t_R _0791_ (.A(net14),
    .Y(_0153_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Right_50 ();
 NAND2x1_ASAP7_75t_R _0793_ (.A(_0153_),
    .B(net15),
    .Y(_0155_));
 OA211x2_ASAP7_75t_R _0794_ (.A1(_0142_),
    .A2(_0152_),
    .B(_0155_),
    .C(net172),
    .Y(_0156_));
 OR3x1_ASAP7_75t_R _0795_ (.A(_0134_),
    .B(_0149_),
    .C(_0156_),
    .Y(_0157_));
 XOR2x1_ASAP7_75t_R _0796_ (.A(net176),
    .Y(_0158_),
    .B(net15));
 NAND3x2_ASAP7_75t_R _0797_ (.B(net10),
    .C(net11),
    .Y(_0159_),
    .A(net176));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Right_49 ();
 NAND2x1_ASAP7_75t_R _0799_ (.A(net2),
    .B(net9),
    .Y(_0161_));
 OR5x1_ASAP7_75t_R _0800_ (.A(net6),
    .B(net2),
    .C(net9),
    .D(net10),
    .E(net11),
    .Y(_0162_));
 OAI21x1_ASAP7_75t_R _0801_ (.A1(_0159_),
    .A2(_0161_),
    .B(_0162_),
    .Y(_0163_));
 NOR2x2_ASAP7_75t_R _0802_ (.A(_0142_),
    .B(_0163_),
    .Y(_0164_));
 XOR2x1_ASAP7_75t_R _0803_ (.A(net6),
    .Y(_0165_),
    .B(net11));
 AND2x2_ASAP7_75t_R _0804_ (.A(_0165_),
    .B(_0133_),
    .Y(_0166_));
 INVx3_ASAP7_75t_R _0805_ (.A(net5),
    .Y(_0167_));
 AND3x1_ASAP7_75t_R _0806_ (.A(_0167_),
    .B(_0146_),
    .C(net4),
    .Y(_0168_));
 AO21x1_ASAP7_75t_R _0807_ (.A1(_0123_),
    .A2(_0132_),
    .B(_0168_),
    .Y(_0169_));
 AOI221x1_ASAP7_75t_R _0808_ (.A1(_0133_),
    .A2(_0158_),
    .B1(_0164_),
    .B2(_0166_),
    .C(_0169_),
    .Y(_0170_));
 AND4x1_ASAP7_75t_R _0809_ (.A(_0122_),
    .B(_0126_),
    .C(_0157_),
    .D(_0170_),
    .Y(_0171_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Right_48 ();
 INVx1_ASAP7_75t_R _0811_ (.A(net9),
    .Y(_0172_));
 INVx2_ASAP7_75t_R _0812_ (.A(net13),
    .Y(_0173_));
 OR4x1_ASAP7_75t_R _0813_ (.A(net172),
    .B(_0173_),
    .C(net14),
    .D(net15),
    .Y(_0174_));
 OAI21x1_ASAP7_75t_R _0814_ (.A1(net13),
    .A2(_0137_),
    .B(_0174_),
    .Y(_0175_));
 AND4x1_ASAP7_75t_R _0815_ (.A(_0146_),
    .B(net9),
    .C(_0150_),
    .D(_0144_),
    .Y(_0176_));
 NOR2x1_ASAP7_75t_R _0816_ (.A(net9),
    .B(_0159_),
    .Y(_0177_));
 OA21x2_ASAP7_75t_R _0817_ (.A1(_0176_),
    .A2(_0177_),
    .B(net97),
    .Y(_0178_));
 AND2x2_ASAP7_75t_R _0818_ (.A(net17),
    .B(_0128_),
    .Y(_0179_));
 AND3x1_ASAP7_75t_R _0819_ (.A(net3),
    .B(net4),
    .C(_0132_),
    .Y(_0180_));
 INVx1_ASAP7_75t_R _0820_ (.A(net17),
    .Y(_0181_));
 AO32x1_ASAP7_75t_R _0821_ (.A1(_0117_),
    .A2(_0123_),
    .A3(_0179_),
    .B1(_0180_),
    .B2(_0181_),
    .Y(_0182_));
 AOI221x1_ASAP7_75t_R _0822_ (.A1(net95),
    .A2(_0175_),
    .B1(_0178_),
    .B2(_0164_),
    .C(_0182_),
    .Y(_0183_));
 AND4x2_ASAP7_75t_R _0823_ (.A(net99),
    .B(net173),
    .C(_0171_),
    .D(_0183_),
    .Y(_0184_));
 AO21x1_ASAP7_75t_R _0824_ (.A1(_0127_),
    .A2(_0130_),
    .B(_0121_),
    .Y(_0185_));
 OAI21x1_ASAP7_75t_R _0825_ (.A1(_0125_),
    .A2(net170),
    .B(_0185_),
    .Y(_0186_));
 AND3x2_ASAP7_75t_R _0826_ (.A(_0171_),
    .B(_0183_),
    .C(_0186_),
    .Y(_0187_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_47 ();
 AO221x1_ASAP7_75t_R _0828_ (.A1(_0172_),
    .A2(_0184_),
    .B1(_0187_),
    .B2(_0173_),
    .C(_0146_),
    .Y(_0189_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_45 ();
 AO221x1_ASAP7_75t_R _0831_ (.A1(net9),
    .A2(_0184_),
    .B1(_0187_),
    .B2(net13),
    .C(net169),
    .Y(_0192_));
 OR3x1_ASAP7_75t_R _0832_ (.A(net2),
    .B(net11),
    .C(_0142_),
    .Y(_0193_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_44 ();
 OR3x1_ASAP7_75t_R _0834_ (.A(net10),
    .B(net13),
    .C(_0153_),
    .Y(_0195_));
 OA211x2_ASAP7_75t_R _0835_ (.A1(net11),
    .A2(net14),
    .B(net15),
    .C(_0195_),
    .Y(_0196_));
 AO21x1_ASAP7_75t_R _0836_ (.A1(net12),
    .A2(_0147_),
    .B(_0196_),
    .Y(_0197_));
 NAND2x1_ASAP7_75t_R _0837_ (.A(_0193_),
    .B(_0197_),
    .Y(_0198_));
 OAI21x1_ASAP7_75t_R _0838_ (.A1(_0137_),
    .A2(_0140_),
    .B(net177),
    .Y(_0199_));
 AND3x1_ASAP7_75t_R _0839_ (.A(net2),
    .B(net11),
    .C(_0199_),
    .Y(_0200_));
 AND3x1_ASAP7_75t_R _0840_ (.A(net10),
    .B(net13),
    .C(_0153_),
    .Y(_0201_));
 AO21x1_ASAP7_75t_R _0841_ (.A1(net11),
    .A2(net14),
    .B(net15),
    .Y(_0202_));
 OA22x2_ASAP7_75t_R _0842_ (.A1(net12),
    .A2(_0147_),
    .B1(_0201_),
    .B2(_0202_),
    .Y(_0203_));
 OR3x1_ASAP7_75t_R _0843_ (.A(net169),
    .B(_0200_),
    .C(_0203_),
    .Y(_0204_));
 OA211x2_ASAP7_75t_R _0844_ (.A1(_0146_),
    .A2(_0198_),
    .B(_0204_),
    .C(net97),
    .Y(_0205_));
 AND3x1_ASAP7_75t_R _0845_ (.A(net169),
    .B(_0127_),
    .C(_0123_),
    .Y(_0206_));
 AO21x1_ASAP7_75t_R _0846_ (.A1(_0146_),
    .A2(net17),
    .B(_0206_),
    .Y(_0207_));
 XOR2x1_ASAP7_75t_R _0847_ (.A(net172),
    .Y(_0208_),
    .B(net14));
 AND3x1_ASAP7_75t_R _0848_ (.A(_0146_),
    .B(net16),
    .C(net4),
    .Y(_0209_));
 AO21x1_ASAP7_75t_R _0849_ (.A1(net172),
    .A2(_0181_),
    .B(_0209_),
    .Y(_0210_));
 AND2x2_ASAP7_75t_R _0850_ (.A(net15),
    .B(_0122_),
    .Y(_0211_));
 AOI21x1_ASAP7_75t_R _0851_ (.A1(_0147_),
    .A2(_0126_),
    .B(_0211_),
    .Y(_0212_));
 AO221x1_ASAP7_75t_R _0852_ (.A1(_0182_),
    .A2(_0208_),
    .B1(_0210_),
    .B2(_0167_),
    .C(_0212_),
    .Y(_0213_));
 AO21x1_ASAP7_75t_R _0853_ (.A1(net5),
    .A2(_0207_),
    .B(_0213_),
    .Y(_0214_));
 AOI211x1_ASAP7_75t_R _0854_ (.A1(_0189_),
    .A2(_0192_),
    .B(_0205_),
    .C(_0214_),
    .Y(_0721_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_42 ();
 NOR2x1_ASAP7_75t_R _0857_ (.A(net24),
    .B(net20),
    .Y(_0217_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_39 ();
 OR3x1_ASAP7_75t_R _0861_ (.A(net32),
    .B(net33),
    .C(net19),
    .Y(_0221_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_38 ();
 AND2x2_ASAP7_75t_R _0863_ (.A(net24),
    .B(net20),
    .Y(_0223_));
 NAND3x1_ASAP7_75t_R _0864_ (.A(net32),
    .B(net33),
    .C(net19),
    .Y(_0224_));
 AO22x1_ASAP7_75t_R _0865_ (.A1(_0217_),
    .A2(_0221_),
    .B1(_0223_),
    .B2(_0224_),
    .Y(_0225_));
 INVx3_ASAP7_75t_R _0866_ (.A(net27),
    .Y(_0226_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_37 ();
 AND5x2_ASAP7_75t_R _0868_ (.A(net24),
    .B(net28),
    .C(net29),
    .D(net30),
    .E(net31),
    .Y(_0228_));
 NAND2x2_ASAP7_75t_R _0869_ (.A(net24),
    .B(net20),
    .Y(_0229_));
 INVx2_ASAP7_75t_R _0870_ (.A(net31),
    .Y(_0230_));
 AOI211x1_ASAP7_75t_R _0871_ (.A1(_0226_),
    .A2(_0228_),
    .B(_0229_),
    .C(_0230_),
    .Y(_0231_));
 OR5x2_ASAP7_75t_R _0872_ (.A(net24),
    .B(net28),
    .C(net29),
    .D(net30),
    .E(net31),
    .Y(_0232_));
 OA211x2_ASAP7_75t_R _0873_ (.A1(_0226_),
    .A2(_0232_),
    .B(_0217_),
    .C(_0230_),
    .Y(_0233_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_36 ();
 NOR2x2_ASAP7_75t_R _0875_ (.A(net21),
    .B(net23),
    .Y(_0235_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_35 ();
 NOR2x1_ASAP7_75t_R _0877_ (.A(net24),
    .B(net22),
    .Y(_0237_));
 AND4x1_ASAP7_75t_R _0878_ (.A(net24),
    .B(net21),
    .C(net22),
    .D(net23),
    .Y(_0238_));
 AOI21x1_ASAP7_75t_R _0879_ (.A1(_0235_),
    .A2(_0237_),
    .B(_0238_),
    .Y(_0239_));
 OR4x2_ASAP7_75t_R _0880_ (.A(_0225_),
    .B(_0231_),
    .C(_0233_),
    .D(_0239_),
    .Y(_0240_));
 INVx6_ASAP7_75t_R _0881_ (.A(net24),
    .Y(_0241_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_34 ();
 OR3x1_ASAP7_75t_R _0883_ (.A(_0241_),
    .B(net26),
    .C(_0226_),
    .Y(_0243_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_33 ();
 INVx1_ASAP7_75t_R _0885_ (.A(net26),
    .Y(_0245_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_32 ();
 OR3x1_ASAP7_75t_R _0887_ (.A(net24),
    .B(_0245_),
    .C(net27),
    .Y(_0247_));
 NAND2x1_ASAP7_75t_R _0888_ (.A(_0243_),
    .B(_0247_),
    .Y(_0248_));
 OR5x1_ASAP7_75t_R _0889_ (.A(net24),
    .B(net32),
    .C(net33),
    .D(net19),
    .E(net20),
    .Y(_0249_));
 OA21x2_ASAP7_75t_R _0890_ (.A1(_0229_),
    .A2(_0224_),
    .B(_0249_),
    .Y(_0250_));
 OR2x6_ASAP7_75t_R _0891_ (.A(_0250_),
    .B(_0239_),
    .Y(_0251_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_31 ();
 INVx8_ASAP7_75t_R _0893_ (.A(_0251_),
    .Y(_0695_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_29 ();
 NOR3x1_ASAP7_75t_R _0896_ (.A(net24),
    .B(net30),
    .C(net31),
    .Y(_0255_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 NOR2x1_ASAP7_75t_R _0898_ (.A(net28),
    .B(net29),
    .Y(_0257_));
 AO21x2_ASAP7_75t_R _0899_ (.A1(_0255_),
    .A2(_0257_),
    .B(_0228_),
    .Y(_0258_));
 AND3x1_ASAP7_75t_R _0900_ (.A(_0248_),
    .B(_0695_),
    .C(_0258_),
    .Y(_0259_));
 INVx1_ASAP7_75t_R _0901_ (.A(_0259_),
    .Y(_0260_));
 INVx1_ASAP7_75t_R _0902_ (.A(net20),
    .Y(_0261_));
 OR3x1_ASAP7_75t_R _0903_ (.A(_0241_),
    .B(net19),
    .C(_0261_),
    .Y(_0262_));
 INVx1_ASAP7_75t_R _0904_ (.A(net19),
    .Y(_0263_));
 OR3x1_ASAP7_75t_R _0905_ (.A(net24),
    .B(_0263_),
    .C(net20),
    .Y(_0264_));
 AO21x1_ASAP7_75t_R _0906_ (.A1(_0262_),
    .A2(_0264_),
    .B(_0239_),
    .Y(_0265_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 XNOR2x1_ASAP7_75t_R _0908_ (.B(net23),
    .Y(_0267_),
    .A(net24));
 OR3x1_ASAP7_75t_R _0909_ (.A(_0241_),
    .B(net30),
    .C(_0230_),
    .Y(_0268_));
 INVx1_ASAP7_75t_R _0910_ (.A(net30),
    .Y(_0269_));
 OR3x1_ASAP7_75t_R _0911_ (.A(net24),
    .B(_0269_),
    .C(net31),
    .Y(_0270_));
 AO21x1_ASAP7_75t_R _0912_ (.A1(_0268_),
    .A2(_0270_),
    .B(_0251_),
    .Y(_0271_));
 AND4x2_ASAP7_75t_R _0913_ (.A(_0260_),
    .B(_0265_),
    .C(_0267_),
    .D(_0271_),
    .Y(_0272_));
 NAND2x1_ASAP7_75t_R _0914_ (.A(_0240_),
    .B(_0272_),
    .Y(_0724_));
 INVx1_ASAP7_75t_R _0915_ (.A(_0724_),
    .Y(_0692_));
 AND2x2_ASAP7_75t_R _0916_ (.A(net28),
    .B(net29),
    .Y(_0273_));
 NOR2x1_ASAP7_75t_R _0917_ (.A(net30),
    .B(net31),
    .Y(_0274_));
 AND2x2_ASAP7_75t_R _0918_ (.A(net30),
    .B(net31),
    .Y(_0275_));
 AO21x1_ASAP7_75t_R _0919_ (.A1(_0273_),
    .A2(_0274_),
    .B(_0275_),
    .Y(_0276_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 INVx2_ASAP7_75t_R _0921_ (.A(net25),
    .Y(_0278_));
 OR3x1_ASAP7_75t_R _0922_ (.A(net24),
    .B(net26),
    .C(net27),
    .Y(_0279_));
 NOR2x1_ASAP7_75t_R _0923_ (.A(_0278_),
    .B(_0279_),
    .Y(_0280_));
 AND4x1_ASAP7_75t_R _0924_ (.A(net24),
    .B(_0278_),
    .C(net26),
    .D(net27),
    .Y(_0281_));
 OAI21x1_ASAP7_75t_R _0925_ (.A1(_0280_),
    .A2(_0281_),
    .B(_0258_),
    .Y(_0282_));
 OR2x2_ASAP7_75t_R _0926_ (.A(_0251_),
    .B(_0282_),
    .Y(_0283_));
 INVx1_ASAP7_75t_R _0927_ (.A(_0283_),
    .Y(_0284_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 AO221x1_ASAP7_75t_R _0930_ (.A1(_0695_),
    .A2(_0276_),
    .B1(_0284_),
    .B2(net18),
    .C(net24),
    .Y(_0287_));
 AO21x1_ASAP7_75t_R _0931_ (.A1(_0275_),
    .A2(_0257_),
    .B(_0274_),
    .Y(_0288_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 AOI21x1_ASAP7_75t_R _0933_ (.A1(_0695_),
    .A2(_0288_),
    .B(_0241_),
    .Y(_0290_));
 OAI21x1_ASAP7_75t_R _0934_ (.A1(net18),
    .A2(_0283_),
    .B(_0290_),
    .Y(_0291_));
 AND2x2_ASAP7_75t_R _0935_ (.A(_0287_),
    .B(_0291_),
    .Y(_0292_));
 AO21x2_ASAP7_75t_R _0936_ (.A1(_0235_),
    .A2(_0237_),
    .B(_0238_),
    .Y(_0293_));
 INVx1_ASAP7_75t_R _0937_ (.A(net33),
    .Y(_0294_));
 OR4x2_ASAP7_75t_R _0938_ (.A(net24),
    .B(_0294_),
    .C(net19),
    .D(net20),
    .Y(_0295_));
 OR3x2_ASAP7_75t_R _0939_ (.A(net33),
    .B(_0263_),
    .C(_0229_),
    .Y(_0296_));
 NAND2x2_ASAP7_75t_R _0940_ (.A(_0295_),
    .B(_0296_),
    .Y(_0297_));
 INVx2_ASAP7_75t_R _0941_ (.A(net29),
    .Y(_0298_));
 AND3x1_ASAP7_75t_R _0942_ (.A(net24),
    .B(_0298_),
    .C(_0275_),
    .Y(_0299_));
 AO21x2_ASAP7_75t_R _0943_ (.A1(net29),
    .A2(_0255_),
    .B(_0299_),
    .Y(_0300_));
 INVx2_ASAP7_75t_R _0944_ (.A(net22),
    .Y(_0301_));
 NOR2x1_ASAP7_75t_R _0945_ (.A(_0301_),
    .B(net23),
    .Y(_0302_));
 AND3x1_ASAP7_75t_R _0946_ (.A(net24),
    .B(_0301_),
    .C(net23),
    .Y(_0303_));
 AO21x1_ASAP7_75t_R _0947_ (.A1(_0241_),
    .A2(_0302_),
    .B(_0303_),
    .Y(_0304_));
 AO221x2_ASAP7_75t_R _0948_ (.A1(_0293_),
    .A2(_0297_),
    .B1(_0300_),
    .B2(_0695_),
    .C(_0304_),
    .Y(_0305_));
 OAI21x1_ASAP7_75t_R _0949_ (.A1(net178),
    .A2(_0282_),
    .B(_0240_),
    .Y(_0306_));
 NOR2x2_ASAP7_75t_R _0950_ (.A(_0305_),
    .B(_0306_),
    .Y(_0307_));
 NOR2x2_ASAP7_75t_R _0951_ (.A(_0251_),
    .B(_0258_),
    .Y(_0308_));
 XOR2x1_ASAP7_75t_R _0952_ (.A(net24),
    .Y(_0309_),
    .B(net27));
 AND2x2_ASAP7_75t_R _0953_ (.A(_0293_),
    .B(_0250_),
    .Y(_0310_));
 AO221x1_ASAP7_75t_R _0954_ (.A1(_0261_),
    .A2(_0239_),
    .B1(_0310_),
    .B2(_0230_),
    .C(_0241_),
    .Y(_0311_));
 AO221x1_ASAP7_75t_R _0955_ (.A1(net20),
    .A2(_0239_),
    .B1(_0310_),
    .B2(net31),
    .C(net24),
    .Y(_0312_));
 AO22x1_ASAP7_75t_R _0956_ (.A1(_0308_),
    .A2(_0309_),
    .B1(_0311_),
    .B2(_0312_),
    .Y(_0313_));
 AND3x1_ASAP7_75t_R _0957_ (.A(_0272_),
    .B(_0307_),
    .C(_0313_),
    .Y(_0314_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 OA21x2_ASAP7_75t_R _0959_ (.A1(_0294_),
    .A2(_0261_),
    .B(_0263_),
    .Y(_0316_));
 OA211x2_ASAP7_75t_R _0960_ (.A1(net33),
    .A2(net20),
    .B(net19),
    .C(_0241_),
    .Y(_0317_));
 AO21x1_ASAP7_75t_R _0961_ (.A1(net24),
    .A2(_0316_),
    .B(_0317_),
    .Y(_0318_));
 AOI21x1_ASAP7_75t_R _0962_ (.A1(_0268_),
    .A2(_0270_),
    .B(net178),
    .Y(_0319_));
 NOR2x1_ASAP7_75t_R _0963_ (.A(_0226_),
    .B(_0232_),
    .Y(_0320_));
 AO21x1_ASAP7_75t_R _0964_ (.A1(_0226_),
    .A2(_0228_),
    .B(_0320_),
    .Y(_0321_));
 NAND2x1_ASAP7_75t_R _0965_ (.A(_0695_),
    .B(_0321_),
    .Y(_0322_));
 INVx1_ASAP7_75t_R _0966_ (.A(_0322_),
    .Y(_0323_));
 AO221x1_ASAP7_75t_R _0967_ (.A1(_0298_),
    .A2(_0319_),
    .B1(_0323_),
    .B2(_0245_),
    .C(_0241_),
    .Y(_0324_));
 AO221x1_ASAP7_75t_R _0968_ (.A1(net29),
    .A2(_0319_),
    .B1(_0323_),
    .B2(net26),
    .C(net24),
    .Y(_0325_));
 NAND2x1_ASAP7_75t_R _0969_ (.A(net21),
    .B(net23),
    .Y(_0326_));
 AO32x1_ASAP7_75t_R _0970_ (.A1(net32),
    .A2(_0235_),
    .A3(_0297_),
    .B1(_0326_),
    .B2(net24),
    .Y(_0327_));
 NOR2x1_ASAP7_75t_R _0971_ (.A(net24),
    .B(_0235_),
    .Y(_0328_));
 INVx1_ASAP7_75t_R _0972_ (.A(net32),
    .Y(_0329_));
 AND4x1_ASAP7_75t_R _0973_ (.A(_0329_),
    .B(net21),
    .C(net23),
    .D(_0297_),
    .Y(_0330_));
 OA21x2_ASAP7_75t_R _0974_ (.A1(_0328_),
    .A2(_0330_),
    .B(net22),
    .Y(_0331_));
 AO21x1_ASAP7_75t_R _0975_ (.A1(_0301_),
    .A2(_0327_),
    .B(_0331_),
    .Y(_0332_));
 AO221x1_ASAP7_75t_R _0976_ (.A1(_0293_),
    .A2(_0318_),
    .B1(_0324_),
    .B2(_0325_),
    .C(_0332_),
    .Y(_0333_));
 NAND2x1_ASAP7_75t_R _0977_ (.A(net25),
    .B(_0290_),
    .Y(_0334_));
 OA211x2_ASAP7_75t_R _0978_ (.A1(net25),
    .A2(_0287_),
    .B(_0334_),
    .C(_0259_),
    .Y(_0335_));
 OR4x2_ASAP7_75t_R _0979_ (.A(_0292_),
    .B(_0314_),
    .C(_0333_),
    .D(_0335_),
    .Y(_0701_));
 AND2x2_ASAP7_75t_R _0980_ (.A(net155),
    .B(net167),
    .Y(_0336_));
 INVx2_ASAP7_75t_R _0981_ (.A(net164),
    .Y(_0337_));
 OA21x2_ASAP7_75t_R _0982_ (.A1(_0001_),
    .A2(_0337_),
    .B(_0000_),
    .Y(_0338_));
 MAJx2_ASAP7_75t_R _0983_ (.A(_0307_),
    .B(_0336_),
    .C(_0338_),
    .Y(_0693_));
 OA21x2_ASAP7_75t_R _0984_ (.A1(_0003_),
    .A2(_0693_),
    .B(_0005_),
    .Y(_0339_));
 OA21x2_ASAP7_75t_R _0985_ (.A1(_0004_),
    .A2(_0339_),
    .B(_0006_),
    .Y(_0696_));
 XNOR2x2_ASAP7_75t_R _0986_ (.A(_0004_),
    .B(net101),
    .Y(_0340_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 NOR2x2_ASAP7_75t_R _0990_ (.A(net81),
    .B(net82),
    .Y(_0344_));
 AND2x4_ASAP7_75t_R _0991_ (.A(_0344_),
    .B(_0340_),
    .Y(_0345_));
 OR3x4_ASAP7_75t_R _0992_ (.A(_0002_),
    .B(_0305_),
    .C(_0306_),
    .Y(_0346_));
 OAI21x1_ASAP7_75t_R _0993_ (.A1(_0305_),
    .A2(_0306_),
    .B(net175),
    .Y(_0347_));
 NAND2x1_ASAP7_75t_R _0994_ (.A(_0346_),
    .B(_0347_),
    .Y(_0348_));
 AND3x1_ASAP7_75t_R _0995_ (.A(_0008_),
    .B(net157),
    .C(net168),
    .Y(_0349_));
 NAND2x2_ASAP7_75t_R _0996_ (.A(net156),
    .B(net168),
    .Y(_0350_));
 AND4x1_ASAP7_75t_R _0997_ (.A(_0008_),
    .B(_0350_),
    .C(_0346_),
    .D(_0347_),
    .Y(_0351_));
 INVx2_ASAP7_75t_R _0998_ (.A(net66),
    .Y(_0352_));
 AOI211x1_ASAP7_75t_R _0999_ (.A1(_0348_),
    .A2(_0349_),
    .B(_0351_),
    .C(_0352_),
    .Y(_0353_));
 NAND2x1_ASAP7_75t_R _1000_ (.A(_0345_),
    .B(_0353_),
    .Y(_0354_));
 AND5x1_ASAP7_75t_R _1001_ (.A(net18),
    .B(net24),
    .C(net25),
    .D(net26),
    .E(net27),
    .Y(_0355_));
 OR3x1_ASAP7_75t_R _1002_ (.A(net18),
    .B(net25),
    .C(_0279_),
    .Y(_0356_));
 INVx1_ASAP7_75t_R _1003_ (.A(_0356_),
    .Y(_0357_));
 OA211x2_ASAP7_75t_R _1004_ (.A1(_0355_),
    .A2(_0357_),
    .B(_0695_),
    .C(_0258_),
    .Y(_0358_));
 AND3x2_ASAP7_75t_R _1005_ (.A(net98),
    .B(_0199_),
    .C(_0163_),
    .Y(_0359_));
 XOR2x1_ASAP7_75t_R _1006_ (.A(net169),
    .Y(_0360_),
    .B(net24));
 OR3x4_ASAP7_75t_R _1007_ (.A(_0358_),
    .B(_0359_),
    .C(_0360_),
    .Y(_0361_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 XNOR2x2_ASAP7_75t_R _1009_ (.A(net169),
    .B(net24),
    .Y(_0363_));
 OR3x4_ASAP7_75t_R _1010_ (.A(_0358_),
    .B(_0359_),
    .C(_0363_),
    .Y(_0364_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 AO21x1_ASAP7_75t_R _1012_ (.A1(_0345_),
    .A2(_0353_),
    .B(_0364_),
    .Y(_0366_));
 OA21x2_ASAP7_75t_R _1013_ (.A1(_0354_),
    .A2(_0361_),
    .B(_0366_),
    .Y(_0703_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 AO21x1_ASAP7_75t_R _1017_ (.A1(net18),
    .A2(net8),
    .B(net7),
    .Y(_0370_));
 OAI21x1_ASAP7_75t_R _1018_ (.A1(net169),
    .A2(net7),
    .B(net18),
    .Y(_0371_));
 INVx2_ASAP7_75t_R _1019_ (.A(net8),
    .Y(_0372_));
 AND3x1_ASAP7_75t_R _1020_ (.A(net18),
    .B(net8),
    .C(net7),
    .Y(_0373_));
 AO221x1_ASAP7_75t_R _1021_ (.A1(net169),
    .A2(_0370_),
    .B1(_0371_),
    .B2(_0372_),
    .C(_0373_),
    .Y(_0704_));
 INVx2_ASAP7_75t_R _1022_ (.A(net79),
    .Y(_0374_));
 AND3x2_ASAP7_75t_R _1023_ (.A(net88),
    .B(_0374_),
    .C(net174),
    .Y(_0375_));
 INVx1_ASAP7_75t_R _1024_ (.A(_0375_),
    .Y(_0376_));
 NAND3x2_ASAP7_75t_R _1025_ (.B(_0346_),
    .C(_0347_),
    .Y(_0377_),
    .A(_0350_));
 AO21x2_ASAP7_75t_R _1026_ (.A1(_0346_),
    .A2(_0347_),
    .B(_0350_),
    .Y(_0378_));
 NAND2x2_ASAP7_75t_R _1027_ (.A(net102),
    .B(_0378_),
    .Y(_0379_));
 INVx2_ASAP7_75t_R _1028_ (.A(_0007_),
    .Y(_0380_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 NAND2x2_ASAP7_75t_R _1030_ (.A(_0380_),
    .B(net70),
    .Y(_0382_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 INVx1_ASAP7_75t_R _1033_ (.A(_0008_),
    .Y(_0385_));
 AND2x2_ASAP7_75t_R _1034_ (.A(net67),
    .B(_0080_),
    .Y(_0386_));
 AO21x2_ASAP7_75t_R _1035_ (.A1(_0385_),
    .A2(_0352_),
    .B(_0386_),
    .Y(_0387_));
 AO21x2_ASAP7_75t_R _1036_ (.A1(net102),
    .A2(net103),
    .B(_0387_),
    .Y(_0388_));
 OAI21x1_ASAP7_75t_R _1037_ (.A1(_0379_),
    .A2(_0382_),
    .B(_0388_),
    .Y(_0389_));
 NOR2x2_ASAP7_75t_R _1038_ (.A(_0358_),
    .B(_0359_),
    .Y(_0390_));
 AND2x6_ASAP7_75t_R _1039_ (.A(_0390_),
    .B(_0360_),
    .Y(_0391_));
 OA21x2_ASAP7_75t_R _1040_ (.A1(_0376_),
    .A2(net94),
    .B(_0391_),
    .Y(_0392_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 NOR3x1_ASAP7_75t_R _1042_ (.A(_0361_),
    .B(_0376_),
    .C(net93),
    .Y(_0394_));
 OR2x2_ASAP7_75t_R _1043_ (.A(_0392_),
    .B(_0394_),
    .Y(_0711_));
 AND2x2_ASAP7_75t_R _1044_ (.A(net88),
    .B(_0374_),
    .Y(_0395_));
 INVx1_ASAP7_75t_R _1045_ (.A(_0395_),
    .Y(_0396_));
 AND2x2_ASAP7_75t_R _1046_ (.A(_0340_),
    .B(_0387_),
    .Y(_0397_));
 XOR2x2_ASAP7_75t_R _1047_ (.A(_0004_),
    .B(net101),
    .Y(_0398_));
 AND3x1_ASAP7_75t_R _1048_ (.A(_0007_),
    .B(_0352_),
    .C(_0340_),
    .Y(_0399_));
 AO221x1_ASAP7_75t_R _1049_ (.A1(net67),
    .A2(_0398_),
    .B1(_0377_),
    .B2(net103),
    .C(_0399_),
    .Y(_0400_));
 OAI21x1_ASAP7_75t_R _1050_ (.A1(_0379_),
    .A2(_0397_),
    .B(_0400_),
    .Y(_0401_));
 OAI21x1_ASAP7_75t_R _1051_ (.A1(_0396_),
    .A2(_0401_),
    .B(_0391_),
    .Y(_0402_));
 OR3x1_ASAP7_75t_R _1052_ (.A(_0361_),
    .B(_0396_),
    .C(_0401_),
    .Y(_0403_));
 NAND2x1_ASAP7_75t_R _1053_ (.A(_0402_),
    .B(_0403_),
    .Y(_0730_));
 AND2x4_ASAP7_75t_R _1054_ (.A(_0390_),
    .B(_0363_),
    .Y(_0404_));
 AO21x2_ASAP7_75t_R _1055_ (.A1(_0377_),
    .A2(net103),
    .B(_0385_),
    .Y(_0405_));
 AND3x2_ASAP7_75t_R _1056_ (.A(net82),
    .B(_0374_),
    .C(_0398_),
    .Y(_0406_));
 AND2x2_ASAP7_75t_R _1057_ (.A(_0007_),
    .B(_0352_),
    .Y(_0407_));
 NAND3x2_ASAP7_75t_R _1058_ (.B(_0378_),
    .C(_0407_),
    .Y(_0408_),
    .A(net102));
 NAND2x1_ASAP7_75t_R _1059_ (.A(_0352_),
    .B(_0080_),
    .Y(_0409_));
 AO21x2_ASAP7_75t_R _1060_ (.A1(_0377_),
    .A2(_0378_),
    .B(_0409_),
    .Y(_0410_));
 NAND2x2_ASAP7_75t_R _1061_ (.A(_0408_),
    .B(_0410_),
    .Y(_0411_));
 AO32x1_ASAP7_75t_R _1062_ (.A1(net75),
    .A2(_0405_),
    .A3(_0406_),
    .B1(_0411_),
    .B2(_0375_),
    .Y(_0412_));
 AOI221x1_ASAP7_75t_R _1063_ (.A1(_0375_),
    .A2(_0411_),
    .B1(_0406_),
    .B2(_0353_),
    .C(_0364_),
    .Y(_0413_));
 AO21x1_ASAP7_75t_R _1064_ (.A1(_0404_),
    .A2(_0412_),
    .B(_0413_),
    .Y(_0728_));
 INVx2_ASAP7_75t_R _1065_ (.A(net82),
    .Y(_0414_));
 OR3x4_ASAP7_75t_R _1066_ (.A(_0414_),
    .B(net77),
    .C(_0340_),
    .Y(_0415_));
 OA21x2_ASAP7_75t_R _1067_ (.A1(net93),
    .A2(_0415_),
    .B(_0391_),
    .Y(_0416_));
 NOR3x2_ASAP7_75t_R _1068_ (.B(net93),
    .C(_0415_),
    .Y(_0417_),
    .A(_0361_));
 OR2x2_ASAP7_75t_R _1069_ (.A(_0416_),
    .B(_0417_),
    .Y(_0734_));
 XOR2x2_ASAP7_75t_R _1070_ (.A(net169),
    .B(net7),
    .Y(_0418_));
 XOR2x1_ASAP7_75t_R _1071_ (.A(net19),
    .Y(_0419_),
    .B(net8));
 AND3x4_ASAP7_75t_R _1072_ (.A(net169),
    .B(_0372_),
    .C(net7),
    .Y(_0420_));
 OR3x4_ASAP7_75t_R _1073_ (.A(net169),
    .B(_0372_),
    .C(net7),
    .Y(_0421_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 NOR2x1_ASAP7_75t_R _1075_ (.A(net33),
    .B(_0421_),
    .Y(_0423_));
 AO221x1_ASAP7_75t_R _1076_ (.A1(_0418_),
    .A2(_0419_),
    .B1(_0420_),
    .B2(net33),
    .C(_0423_),
    .Y(_0735_));
 INVx1_ASAP7_75t_R _1077_ (.A(_0735_),
    .Y(_0715_));
 AND3x1_ASAP7_75t_R _1078_ (.A(net76),
    .B(net77),
    .C(net174),
    .Y(_0424_));
 AND3x1_ASAP7_75t_R _1079_ (.A(_0374_),
    .B(_0398_),
    .C(_0407_),
    .Y(_0425_));
 NOR2x1_ASAP7_75t_R _1080_ (.A(_0424_),
    .B(_0425_),
    .Y(_0426_));
 NOR2x1_ASAP7_75t_R _1081_ (.A(_0414_),
    .B(_0426_),
    .Y(_0427_));
 AND4x1_ASAP7_75t_R _1082_ (.A(net102),
    .B(net103),
    .C(_0387_),
    .D(_0406_),
    .Y(_0428_));
 AO21x1_ASAP7_75t_R _1083_ (.A1(_0379_),
    .A2(_0427_),
    .B(_0428_),
    .Y(_0429_));
 NAND2x1_ASAP7_75t_R _1084_ (.A(_0404_),
    .B(_0429_),
    .Y(_0430_));
 OAI21x1_ASAP7_75t_R _1085_ (.A1(_0364_),
    .A2(_0429_),
    .B(_0430_),
    .Y(_0738_));
 AO21x1_ASAP7_75t_R _1086_ (.A1(_0408_),
    .A2(_0410_),
    .B(_0415_),
    .Y(_0431_));
 AND2x2_ASAP7_75t_R _1087_ (.A(net85),
    .B(net79),
    .Y(_0432_));
 AND2x4_ASAP7_75t_R _1088_ (.A(_0340_),
    .B(_0432_),
    .Y(_0433_));
 NAND2x1_ASAP7_75t_R _1089_ (.A(_0353_),
    .B(_0433_),
    .Y(_0434_));
 NAND2x1_ASAP7_75t_R _1090_ (.A(_0431_),
    .B(_0434_),
    .Y(_0435_));
 AND3x1_ASAP7_75t_R _1091_ (.A(_0391_),
    .B(_0431_),
    .C(_0434_),
    .Y(_0436_));
 AO21x1_ASAP7_75t_R _1092_ (.A1(_0404_),
    .A2(_0435_),
    .B(_0436_),
    .Y(_0736_));
 INVx2_ASAP7_75t_R _1093_ (.A(_0433_),
    .Y(_0437_));
 OA21x2_ASAP7_75t_R _1094_ (.A1(net93),
    .A2(_0437_),
    .B(_0391_),
    .Y(_0438_));
 NOR3x2_ASAP7_75t_R _1095_ (.B(net93),
    .C(_0437_),
    .Y(_0439_),
    .A(_0361_));
 OR2x2_ASAP7_75t_R _1096_ (.A(_0438_),
    .B(_0439_),
    .Y(_0742_));
 XOR2x1_ASAP7_75t_R _1097_ (.A(net30),
    .Y(_0440_),
    .B(net8));
 NOR2x1_ASAP7_75t_R _1098_ (.A(net29),
    .B(_0421_),
    .Y(_0441_));
 AO221x1_ASAP7_75t_R _1099_ (.A1(net29),
    .A2(_0420_),
    .B1(_0440_),
    .B2(_0418_),
    .C(_0441_),
    .Y(_0743_));
 INVx1_ASAP7_75t_R _1100_ (.A(_0743_),
    .Y(_0717_));
 NAND2x1_ASAP7_75t_R _1101_ (.A(net86),
    .B(net80),
    .Y(_0442_));
 OAI21x1_ASAP7_75t_R _1102_ (.A1(_0401_),
    .A2(_0442_),
    .B(_0391_),
    .Y(_0443_));
 OR3x1_ASAP7_75t_R _1103_ (.A(_0361_),
    .B(_0401_),
    .C(_0442_),
    .Y(_0444_));
 NAND2x1_ASAP7_75t_R _1104_ (.A(_0443_),
    .B(_0444_),
    .Y(_0746_));
 AND2x4_ASAP7_75t_R _1105_ (.A(_0398_),
    .B(_0432_),
    .Y(_0445_));
 AO32x1_ASAP7_75t_R _1106_ (.A1(net74),
    .A2(_0405_),
    .A3(_0445_),
    .B1(_0433_),
    .B2(_0411_),
    .Y(_0446_));
 AOI221x1_ASAP7_75t_R _1107_ (.A1(_0411_),
    .A2(_0433_),
    .B1(_0445_),
    .B2(_0353_),
    .C(_0364_),
    .Y(_0447_));
 AO21x1_ASAP7_75t_R _1108_ (.A1(_0404_),
    .A2(_0446_),
    .B(_0447_),
    .Y(_0744_));
 OR2x2_ASAP7_75t_R _1109_ (.A(_0025_),
    .B(_0083_),
    .Y(_0448_));
 OA21x2_ASAP7_75t_R _1110_ (.A1(_0027_),
    .A2(_0028_),
    .B(_0026_),
    .Y(_0449_));
 OR5x1_ASAP7_75t_R _1111_ (.A(_0025_),
    .B(_0027_),
    .C(_0029_),
    .D(_0030_),
    .E(_0083_),
    .Y(_0450_));
 OA211x2_ASAP7_75t_R _1112_ (.A1(_0448_),
    .A2(_0449_),
    .B(_0450_),
    .C(_0024_),
    .Y(_0451_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 OR2x2_ASAP7_75t_R _1114_ (.A(_0021_),
    .B(_0023_),
    .Y(_0452_));
 OA21x2_ASAP7_75t_R _1115_ (.A1(_0021_),
    .A2(_0022_),
    .B(_0020_),
    .Y(_0453_));
 OA21x2_ASAP7_75t_R _1116_ (.A1(_0451_),
    .A2(_0452_),
    .B(_0453_),
    .Y(_0454_));
 OR3x1_ASAP7_75t_R _1117_ (.A(_0019_),
    .B(_0082_),
    .C(_0454_),
    .Y(_0455_));
 AND2x2_ASAP7_75t_R _1118_ (.A(_0018_),
    .B(_0455_),
    .Y(_0713_));
 OR4x1_ASAP7_75t_R _1119_ (.A(_0015_),
    .B(_0017_),
    .C(_0019_),
    .D(_0082_),
    .Y(_0456_));
 OA21x2_ASAP7_75t_R _1120_ (.A1(_0017_),
    .A2(_0018_),
    .B(_0016_),
    .Y(_0457_));
 OA21x2_ASAP7_75t_R _1121_ (.A1(_0015_),
    .A2(_0457_),
    .B(_0014_),
    .Y(_0458_));
 OA21x2_ASAP7_75t_R _1122_ (.A1(_0454_),
    .A2(_0456_),
    .B(_0458_),
    .Y(_0459_));
 OR3x1_ASAP7_75t_R _1123_ (.A(_0013_),
    .B(_0012_),
    .C(_0459_),
    .Y(_0460_));
 NAND2x1_ASAP7_75t_R _1124_ (.A(_0460_),
    .B(_0011_),
    .Y(_0710_));
 INVx1_ASAP7_75t_R _1125_ (.A(_0040_),
    .Y(net58));
 INVx1_ASAP7_75t_R _1126_ (.A(_0041_),
    .Y(net57));
 INVx1_ASAP7_75t_R _1127_ (.A(_0042_),
    .Y(net55));
 INVx1_ASAP7_75t_R _1128_ (.A(_0043_),
    .Y(net54));
 INVx1_ASAP7_75t_R _1129_ (.A(_0044_),
    .Y(net53));
 INVx1_ASAP7_75t_R _1130_ (.A(_0045_),
    .Y(net52));
 INVx1_ASAP7_75t_R _1131_ (.A(_0046_),
    .Y(net51));
 INVx1_ASAP7_75t_R _1132_ (.A(_0047_),
    .Y(net50));
 INVx1_ASAP7_75t_R _1133_ (.A(_0048_),
    .Y(net49));
 INVx1_ASAP7_75t_R _1134_ (.A(_0049_),
    .Y(net48));
 INVx1_ASAP7_75t_R _1135_ (.A(_0050_),
    .Y(net47));
 INVx1_ASAP7_75t_R _1136_ (.A(_0051_),
    .Y(net46));
 INVx1_ASAP7_75t_R _1137_ (.A(_0052_),
    .Y(net44));
 INVx1_ASAP7_75t_R _1138_ (.A(_0053_),
    .Y(net43));
 INVx1_ASAP7_75t_R _1139_ (.A(_0054_),
    .Y(net42));
 INVx1_ASAP7_75t_R _1140_ (.A(_0055_),
    .Y(net41));
 INVx1_ASAP7_75t_R _1141_ (.A(_0056_),
    .Y(net40));
 INVx1_ASAP7_75t_R _1142_ (.A(_0057_),
    .Y(net39));
 INVx1_ASAP7_75t_R _1143_ (.A(_0058_),
    .Y(net38));
 INVx1_ASAP7_75t_R _1144_ (.A(_0059_),
    .Y(net37));
 INVx1_ASAP7_75t_R _1145_ (.A(_0060_),
    .Y(net36));
 INVx1_ASAP7_75t_R _1146_ (.A(_0061_),
    .Y(net35));
 INVx1_ASAP7_75t_R _1147_ (.A(_0062_),
    .Y(net65));
 INVx1_ASAP7_75t_R _1148_ (.A(_0063_),
    .Y(net64));
 INVx1_ASAP7_75t_R _1149_ (.A(_0064_),
    .Y(net63));
 INVx1_ASAP7_75t_R _1150_ (.A(_0065_),
    .Y(net62));
 INVx1_ASAP7_75t_R _1151_ (.A(_0066_),
    .Y(net61));
 INVx1_ASAP7_75t_R _1152_ (.A(_0067_),
    .Y(net60));
 INVx1_ASAP7_75t_R _1153_ (.A(_0068_),
    .Y(net59));
 INVx1_ASAP7_75t_R _1154_ (.A(_0069_),
    .Y(net56));
 INVx1_ASAP7_75t_R _1155_ (.A(_0070_),
    .Y(net45));
 INVx1_ASAP7_75t_R _1156_ (.A(_0071_),
    .Y(net34));
 NOR2x1_ASAP7_75t_R _1157_ (.A(_0438_),
    .B(_0439_),
    .Y(_0716_));
 XOR2x1_ASAP7_75t_R _1158_ (.A(net24),
    .Y(_0461_),
    .B(net26));
 AO221x1_ASAP7_75t_R _1159_ (.A1(_0263_),
    .A2(_0239_),
    .B1(_0310_),
    .B2(_0269_),
    .C(_0241_),
    .Y(_0462_));
 AO221x1_ASAP7_75t_R _1160_ (.A1(net19),
    .A2(_0239_),
    .B1(_0310_),
    .B2(net30),
    .C(net24),
    .Y(_0463_));
 AO22x1_ASAP7_75t_R _1161_ (.A1(_0308_),
    .A2(_0461_),
    .B1(_0462_),
    .B2(_0463_),
    .Y(_0464_));
 INVx1_ASAP7_75t_R _1162_ (.A(_0265_),
    .Y(_0465_));
 AO21x2_ASAP7_75t_R _1163_ (.A1(_0295_),
    .A2(_0296_),
    .B(_0239_),
    .Y(_0466_));
 OAI21x1_ASAP7_75t_R _1164_ (.A1(_0298_),
    .A2(net178),
    .B(_0466_),
    .Y(_0467_));
 AND3x1_ASAP7_75t_R _1165_ (.A(_0248_),
    .B(_0695_),
    .C(_0258_),
    .Y(_0468_));
 AO221x1_ASAP7_75t_R _1166_ (.A1(net28),
    .A2(_0319_),
    .B1(_0468_),
    .B2(net18),
    .C(net24),
    .Y(_0469_));
 AO221x1_ASAP7_75t_R _1167_ (.A1(net32),
    .A2(_0465_),
    .B1(_0467_),
    .B2(net31),
    .C(_0469_),
    .Y(_0470_));
 NOR2x1_ASAP7_75t_R _1168_ (.A(net28),
    .B(_0271_),
    .Y(_0471_));
 OAI21x1_ASAP7_75t_R _1169_ (.A1(net29),
    .A2(net178),
    .B(_0466_),
    .Y(_0472_));
 AO22x1_ASAP7_75t_R _1170_ (.A1(_0329_),
    .A2(_0465_),
    .B1(_0472_),
    .B2(_0230_),
    .Y(_0473_));
 INVx1_ASAP7_75t_R _1171_ (.A(net18),
    .Y(_0474_));
 AND2x2_ASAP7_75t_R _1172_ (.A(_0474_),
    .B(_0468_),
    .Y(_0475_));
 OR4x1_ASAP7_75t_R _1173_ (.A(_0241_),
    .B(_0471_),
    .C(_0473_),
    .D(_0475_),
    .Y(_0476_));
 AO32x1_ASAP7_75t_R _1174_ (.A1(_0272_),
    .A2(_0307_),
    .A3(_0464_),
    .B1(_0470_),
    .B2(_0476_),
    .Y(_0477_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 OR3x1_ASAP7_75t_R _1176_ (.A(net33),
    .B(net20),
    .C(_0326_),
    .Y(_0479_));
 INVx1_ASAP7_75t_R _1177_ (.A(_0479_),
    .Y(_0480_));
 AND3x1_ASAP7_75t_R _1178_ (.A(net33),
    .B(net20),
    .C(_0235_),
    .Y(_0481_));
 NAND2x1_ASAP7_75t_R _1179_ (.A(_0301_),
    .B(net23),
    .Y(_0482_));
 OAI22x1_ASAP7_75t_R _1180_ (.A1(net21),
    .A2(net23),
    .B1(_0482_),
    .B2(net20),
    .Y(_0483_));
 AO221x1_ASAP7_75t_R _1181_ (.A1(net21),
    .A2(net23),
    .B1(_0302_),
    .B2(net20),
    .C(net24),
    .Y(_0484_));
 OA21x2_ASAP7_75t_R _1182_ (.A1(_0241_),
    .A2(_0483_),
    .B(_0484_),
    .Y(_0485_));
 AO221x1_ASAP7_75t_R _1183_ (.A1(_0226_),
    .A2(_0300_),
    .B1(_0321_),
    .B2(_0278_),
    .C(_0241_),
    .Y(_0486_));
 AO221x1_ASAP7_75t_R _1184_ (.A1(net27),
    .A2(_0300_),
    .B1(_0321_),
    .B2(net25),
    .C(net24),
    .Y(_0487_));
 AND3x1_ASAP7_75t_R _1185_ (.A(_0695_),
    .B(_0486_),
    .C(_0487_),
    .Y(_0488_));
 OR4x2_ASAP7_75t_R _1186_ (.A(_0480_),
    .B(_0481_),
    .C(_0485_),
    .D(_0488_),
    .Y(_0489_));
 NOR2x2_ASAP7_75t_R _1187_ (.A(_0477_),
    .B(_0489_),
    .Y(_0698_));
 NOR2x1_ASAP7_75t_R _1188_ (.A(_0416_),
    .B(_0417_),
    .Y(_0714_));
 AND4x1_ASAP7_75t_R _1189_ (.A(_0167_),
    .B(net16),
    .C(net3),
    .D(_0123_),
    .Y(_0490_));
 AND3x1_ASAP7_75t_R _1190_ (.A(net13),
    .B(net15),
    .C(net96),
    .Y(_0491_));
 OR3x1_ASAP7_75t_R _1191_ (.A(net172),
    .B(_0490_),
    .C(_0491_),
    .Y(_0492_));
 AO21x1_ASAP7_75t_R _1192_ (.A1(net10),
    .A2(_0184_),
    .B(_0492_),
    .Y(_0493_));
 OR4x1_ASAP7_75t_R _1193_ (.A(_0167_),
    .B(net16),
    .C(net3),
    .D(_0123_),
    .Y(_0494_));
 OR3x1_ASAP7_75t_R _1194_ (.A(net13),
    .B(net15),
    .C(_0134_),
    .Y(_0495_));
 AND3x1_ASAP7_75t_R _1195_ (.A(net169),
    .B(_0494_),
    .C(_0495_),
    .Y(_0496_));
 NAND2x1_ASAP7_75t_R _1196_ (.A(net14),
    .B(_0496_),
    .Y(_0497_));
 AO21x1_ASAP7_75t_R _1197_ (.A1(_0150_),
    .A2(_0184_),
    .B(_0497_),
    .Y(_0498_));
 OA211x2_ASAP7_75t_R _1198_ (.A1(net14),
    .A2(_0493_),
    .B(_0498_),
    .C(_0187_),
    .Y(_0499_));
 INVx1_ASAP7_75t_R _1199_ (.A(net2),
    .Y(_0500_));
 NAND2x1_ASAP7_75t_R _1200_ (.A(net9),
    .B(net11),
    .Y(_0501_));
 OAI21x1_ASAP7_75t_R _1201_ (.A1(_0500_),
    .A2(_0145_),
    .B(_0501_),
    .Y(_0502_));
 OR2x2_ASAP7_75t_R _1202_ (.A(net9),
    .B(net11),
    .Y(_0503_));
 OA211x2_ASAP7_75t_R _1203_ (.A1(net2),
    .A2(_0152_),
    .B(_0503_),
    .C(net172),
    .Y(_0504_));
 INVx1_ASAP7_75t_R _1204_ (.A(_0504_),
    .Y(_0505_));
 OA211x2_ASAP7_75t_R _1205_ (.A1(net169),
    .A2(_0502_),
    .B(_0505_),
    .C(_0199_),
    .Y(_0506_));
 NOR2x1_ASAP7_75t_R _1206_ (.A(net12),
    .B(net14),
    .Y(_0507_));
 AND3x1_ASAP7_75t_R _1207_ (.A(_0144_),
    .B(_0173_),
    .C(net14),
    .Y(_0508_));
 OA211x2_ASAP7_75t_R _1208_ (.A1(_0507_),
    .A2(_0508_),
    .B(net169),
    .C(net15),
    .Y(_0509_));
 AND3x1_ASAP7_75t_R _1209_ (.A(net11),
    .B(net13),
    .C(_0153_),
    .Y(_0510_));
 AO21x1_ASAP7_75t_R _1210_ (.A1(net12),
    .A2(net14),
    .B(_0510_),
    .Y(_0511_));
 AND3x1_ASAP7_75t_R _1211_ (.A(_0146_),
    .B(_0147_),
    .C(_0511_),
    .Y(_0512_));
 OR3x1_ASAP7_75t_R _1212_ (.A(_0506_),
    .B(_0509_),
    .C(_0512_),
    .Y(_0513_));
 INVx1_ASAP7_75t_R _1213_ (.A(_0496_),
    .Y(_0514_));
 AND2x2_ASAP7_75t_R _1214_ (.A(_0150_),
    .B(_0492_),
    .Y(_0515_));
 AO21x1_ASAP7_75t_R _1215_ (.A1(net10),
    .A2(_0514_),
    .B(_0515_),
    .Y(_0516_));
 OR2x2_ASAP7_75t_R _1216_ (.A(net17),
    .B(net4),
    .Y(_0517_));
 NOR2x1_ASAP7_75t_R _1217_ (.A(_0167_),
    .B(_0517_),
    .Y(_0518_));
 AO21x1_ASAP7_75t_R _1218_ (.A1(_0167_),
    .A2(_0117_),
    .B(_0518_),
    .Y(_0519_));
 AO22x1_ASAP7_75t_R _1219_ (.A1(net15),
    .A2(_0117_),
    .B1(net4),
    .B2(_0146_),
    .Y(_0520_));
 AO21x1_ASAP7_75t_R _1220_ (.A1(_0147_),
    .A2(_0181_),
    .B(_0146_),
    .Y(_0521_));
 AND2x2_ASAP7_75t_R _1221_ (.A(net5),
    .B(net3),
    .Y(_0522_));
 AO32x1_ASAP7_75t_R _1222_ (.A1(_0167_),
    .A2(net17),
    .A3(_0520_),
    .B1(_0521_),
    .B2(_0522_),
    .Y(_0523_));
 AO221x1_ASAP7_75t_R _1223_ (.A1(_0492_),
    .A2(_0514_),
    .B1(_0519_),
    .B2(net169),
    .C(_0523_),
    .Y(_0524_));
 AO221x1_ASAP7_75t_R _1224_ (.A1(net97),
    .A2(_0513_),
    .B1(_0516_),
    .B2(_0184_),
    .C(_0524_),
    .Y(_0525_));
 NOR2x1_ASAP7_75t_R _1225_ (.A(_0499_),
    .B(_0525_),
    .Y(_0699_));
 AO21x1_ASAP7_75t_R _1226_ (.A1(net169),
    .A2(net7),
    .B(_0372_),
    .Y(_0705_));
 INVx1_ASAP7_75t_R _1227_ (.A(net165),
    .Y(_0723_));
 AO22x1_ASAP7_75t_R _1228_ (.A1(_0121_),
    .A2(_0125_),
    .B1(_0133_),
    .B2(net173),
    .Y(_0725_));
 AND3x1_ASAP7_75t_R _1229_ (.A(net74),
    .B(_0345_),
    .C(_0379_),
    .Y(_0526_));
 XNOR2x1_ASAP7_75t_R _1230_ (.B(_0526_),
    .Y(_0527_),
    .A(_0363_));
 AND2x2_ASAP7_75t_R _1231_ (.A(_0390_),
    .B(_0527_),
    .Y(_0706_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 XOR2x1_ASAP7_75t_R _1233_ (.A(net20),
    .Y(_0529_),
    .B(net8));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 NOR2x1_ASAP7_75t_R _1236_ (.A(net19),
    .B(_0421_),
    .Y(_0532_));
 AO221x1_ASAP7_75t_R _1237_ (.A1(net19),
    .A2(_0420_),
    .B1(_0529_),
    .B2(_0418_),
    .C(_0532_),
    .Y(_0732_));
 AND4x1_ASAP7_75t_R _1238_ (.A(_0385_),
    .B(net68),
    .C(_0377_),
    .D(_0378_),
    .Y(_0533_));
 AOI22x1_ASAP7_75t_R _1239_ (.A1(_0380_),
    .A2(net69),
    .B1(net102),
    .B2(_0378_),
    .Y(_0534_));
 OR2x6_ASAP7_75t_R _1240_ (.A(_0533_),
    .B(_0534_),
    .Y(_0535_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 AND2x2_ASAP7_75t_R _1242_ (.A(_0352_),
    .B(_0080_),
    .Y(_0537_));
 AND3x2_ASAP7_75t_R _1243_ (.A(net102),
    .B(net103),
    .C(_0537_),
    .Y(_0538_));
 AOI22x1_ASAP7_75t_R _1244_ (.A1(_0433_),
    .A2(_0535_),
    .B1(_0538_),
    .B2(_0406_),
    .Y(_0539_));
 AO221x1_ASAP7_75t_R _1245_ (.A1(_0433_),
    .A2(_0535_),
    .B1(_0538_),
    .B2(_0406_),
    .C(_0364_),
    .Y(_0540_));
 OAI21x1_ASAP7_75t_R _1246_ (.A1(_0361_),
    .A2(_0539_),
    .B(_0540_),
    .Y(_0740_));
 AO31x2_ASAP7_75t_R _1247_ (.A1(net102),
    .A2(_0378_),
    .A3(_0537_),
    .B(_0398_),
    .Y(_0541_));
 OA31x2_ASAP7_75t_R _1248_ (.A1(_0340_),
    .A2(_0533_),
    .A3(_0534_),
    .B1(_0541_),
    .Y(_0542_));
 NAND2x1_ASAP7_75t_R _1249_ (.A(_0432_),
    .B(_0542_),
    .Y(_0543_));
 AND3x1_ASAP7_75t_R _1250_ (.A(_0404_),
    .B(_0432_),
    .C(_0542_),
    .Y(_0544_));
 AO21x1_ASAP7_75t_R _1251_ (.A1(_0391_),
    .A2(_0543_),
    .B(_0544_),
    .Y(_0748_));
 INVx1_ASAP7_75t_R _1252_ (.A(_0445_),
    .Y(_0545_));
 NOR2x1_ASAP7_75t_R _1253_ (.A(_0389_),
    .B(_0545_),
    .Y(_0546_));
 OA21x2_ASAP7_75t_R _1254_ (.A1(_0389_),
    .A2(_0545_),
    .B(_0391_),
    .Y(_0547_));
 AO21x1_ASAP7_75t_R _1255_ (.A1(_0404_),
    .A2(_0546_),
    .B(_0547_),
    .Y(_0719_));
 NAND2x1_ASAP7_75t_R _1256_ (.A(_0375_),
    .B(_0535_),
    .Y(_0548_));
 AND3x1_ASAP7_75t_R _1257_ (.A(_0404_),
    .B(_0375_),
    .C(_0535_),
    .Y(_0549_));
 AO21x1_ASAP7_75t_R _1258_ (.A1(_0391_),
    .A2(_0548_),
    .B(_0549_),
    .Y(_0750_));
 AND2x2_ASAP7_75t_R _1259_ (.A(_0272_),
    .B(_0307_),
    .Y(_0550_));
 AO32x1_ASAP7_75t_R _1260_ (.A1(_0298_),
    .A2(_0293_),
    .A3(_0250_),
    .B1(_0308_),
    .B2(_0278_),
    .Y(_0551_));
 XOR2x1_ASAP7_75t_R _1261_ (.A(net24),
    .Y(_0552_),
    .B(net33));
 AO32x1_ASAP7_75t_R _1262_ (.A1(net29),
    .A2(_0293_),
    .A3(_0250_),
    .B1(_0308_),
    .B2(net25),
    .Y(_0553_));
 AND2x2_ASAP7_75t_R _1263_ (.A(_0241_),
    .B(_0553_),
    .Y(_0554_));
 AO221x1_ASAP7_75t_R _1264_ (.A1(net24),
    .A2(_0551_),
    .B1(_0552_),
    .B2(_0239_),
    .C(_0554_),
    .Y(_0555_));
 AO221x1_ASAP7_75t_R _1265_ (.A1(net20),
    .A2(net23),
    .B1(_0302_),
    .B2(net19),
    .C(net24),
    .Y(_0556_));
 OA21x2_ASAP7_75t_R _1266_ (.A1(net28),
    .A2(_0251_),
    .B(_0265_),
    .Y(_0557_));
 OA222x2_ASAP7_75t_R _1267_ (.A1(net20),
    .A2(net23),
    .B1(_0482_),
    .B2(net19),
    .C1(net31),
    .C2(_0557_),
    .Y(_0558_));
 NAND2x1_ASAP7_75t_R _1268_ (.A(net24),
    .B(_0558_),
    .Y(_0559_));
 AO221x1_ASAP7_75t_R _1269_ (.A1(_0226_),
    .A2(_0319_),
    .B1(_0323_),
    .B2(_0474_),
    .C(_0241_),
    .Y(_0560_));
 AO221x1_ASAP7_75t_R _1270_ (.A1(net27),
    .A2(_0319_),
    .B1(_0323_),
    .B2(net18),
    .C(net24),
    .Y(_0561_));
 AO221x1_ASAP7_75t_R _1271_ (.A1(_0329_),
    .A2(_0261_),
    .B1(_0297_),
    .B2(_0269_),
    .C(_0241_),
    .Y(_0562_));
 AO221x1_ASAP7_75t_R _1272_ (.A1(net32),
    .A2(net20),
    .B1(_0297_),
    .B2(net30),
    .C(net24),
    .Y(_0563_));
 AND3x1_ASAP7_75t_R _1273_ (.A(_0293_),
    .B(_0562_),
    .C(_0563_),
    .Y(_0564_));
 AO221x1_ASAP7_75t_R _1274_ (.A1(_0556_),
    .A2(_0559_),
    .B1(_0560_),
    .B2(_0561_),
    .C(_0564_),
    .Y(_0565_));
 AO21x1_ASAP7_75t_R _1275_ (.A1(net28),
    .A2(_0695_),
    .B(_0465_),
    .Y(_0566_));
 AO32x1_ASAP7_75t_R _1276_ (.A1(net26),
    .A2(_0300_),
    .A3(_0308_),
    .B1(_0566_),
    .B2(net31),
    .Y(_0567_));
 AND4x1_ASAP7_75t_R _1277_ (.A(net24),
    .B(_0245_),
    .C(_0300_),
    .D(_0308_),
    .Y(_0568_));
 AO21x1_ASAP7_75t_R _1278_ (.A1(_0241_),
    .A2(_0567_),
    .B(_0568_),
    .Y(_0569_));
 AOI211x1_ASAP7_75t_R _1279_ (.A1(_0550_),
    .A2(_0555_),
    .B(_0565_),
    .C(_0569_),
    .Y(_0722_));
 OR3x1_ASAP7_75t_R _1280_ (.A(net5),
    .B(net16),
    .C(net3),
    .Y(_0570_));
 AO21x1_ASAP7_75t_R _1281_ (.A1(_0517_),
    .A2(_0570_),
    .B(net169),
    .Y(_0571_));
 NAND2x1_ASAP7_75t_R _1282_ (.A(net169),
    .B(net17),
    .Y(_0572_));
 AO21x1_ASAP7_75t_R _1283_ (.A1(_0146_),
    .A2(net3),
    .B(net5),
    .Y(_0573_));
 AO21x1_ASAP7_75t_R _1284_ (.A1(_0572_),
    .A2(_0573_),
    .B(_0123_),
    .Y(_0574_));
 AO21x1_ASAP7_75t_R _1285_ (.A1(net169),
    .A2(net16),
    .B(_0123_),
    .Y(_0575_));
 OA211x2_ASAP7_75t_R _1286_ (.A1(_0146_),
    .A2(net3),
    .B(_0575_),
    .C(net5),
    .Y(_0576_));
 INVx1_ASAP7_75t_R _1287_ (.A(_0576_),
    .Y(_0577_));
 AO21x1_ASAP7_75t_R _1288_ (.A1(net12),
    .A2(_0147_),
    .B(net14),
    .Y(_0578_));
 AO21x1_ASAP7_75t_R _1289_ (.A1(_0500_),
    .A2(net11),
    .B(_0150_),
    .Y(_0579_));
 AND2x2_ASAP7_75t_R _1290_ (.A(_0146_),
    .B(_0503_),
    .Y(_0580_));
 AO21x1_ASAP7_75t_R _1291_ (.A1(net2),
    .A2(_0144_),
    .B(net10),
    .Y(_0581_));
 AO32x1_ASAP7_75t_R _1292_ (.A1(net172),
    .A2(_0501_),
    .A3(_0579_),
    .B1(_0580_),
    .B2(_0581_),
    .Y(_0582_));
 AND4x1_ASAP7_75t_R _1293_ (.A(net12),
    .B(net14),
    .C(net15),
    .D(_0582_),
    .Y(_0583_));
 AO21x1_ASAP7_75t_R _1294_ (.A1(_0146_),
    .A2(_0578_),
    .B(_0583_),
    .Y(_0584_));
 AO21x1_ASAP7_75t_R _1295_ (.A1(_0153_),
    .A2(_0147_),
    .B(_0146_),
    .Y(_0585_));
 AO21x1_ASAP7_75t_R _1296_ (.A1(net14),
    .A2(net15),
    .B(net172),
    .Y(_0586_));
 OAI21x1_ASAP7_75t_R _1297_ (.A1(net12),
    .A2(_0147_),
    .B(net14),
    .Y(_0587_));
 AO32x1_ASAP7_75t_R _1298_ (.A1(_0147_),
    .A2(_0507_),
    .A3(_0582_),
    .B1(_0587_),
    .B2(net172),
    .Y(_0588_));
 AO22x1_ASAP7_75t_R _1299_ (.A1(_0585_),
    .A2(_0586_),
    .B1(_0588_),
    .B2(_0173_),
    .Y(_0589_));
 AO21x1_ASAP7_75t_R _1300_ (.A1(net13),
    .A2(_0584_),
    .B(_0589_),
    .Y(_0590_));
 AO32x1_ASAP7_75t_R _1301_ (.A1(_0571_),
    .A2(_0574_),
    .A3(_0577_),
    .B1(_0590_),
    .B2(_0133_),
    .Y(_0591_));
 AO221x2_ASAP7_75t_R _1302_ (.A1(_0165_),
    .A2(_0184_),
    .B1(_0187_),
    .B2(_0158_),
    .C(_0591_),
    .Y(_0702_));
 OAI21x1_ASAP7_75t_R _1303_ (.A1(_0250_),
    .A2(_0258_),
    .B(_0293_),
    .Y(_0726_));
 XOR2x1_ASAP7_75t_R _1304_ (.A(net25),
    .Y(_0592_),
    .B(net8));
 NOR2x1_ASAP7_75t_R _1305_ (.A(net18),
    .B(_0421_),
    .Y(_0593_));
 AO221x1_ASAP7_75t_R _1306_ (.A1(net18),
    .A2(_0420_),
    .B1(_0592_),
    .B2(_0418_),
    .C(_0593_),
    .Y(_0707_));
 XOR2x1_ASAP7_75t_R _1307_ (.A(net23),
    .Y(_0594_),
    .B(net8));
 NOR2x1_ASAP7_75t_R _1308_ (.A(net22),
    .B(_0421_),
    .Y(_0595_));
 AO221x2_ASAP7_75t_R _1309_ (.A1(net22),
    .A2(_0420_),
    .B1(_0594_),
    .B2(_0418_),
    .C(_0595_),
    .Y(_0712_));
 XOR2x1_ASAP7_75t_R _1310_ (.A(net21),
    .Y(_0596_),
    .B(net8));
 NOR2x1_ASAP7_75t_R _1311_ (.A(net20),
    .B(_0421_),
    .Y(_0597_));
 AO221x1_ASAP7_75t_R _1312_ (.A1(net20),
    .A2(_0420_),
    .B1(_0596_),
    .B2(_0418_),
    .C(_0597_),
    .Y(_0729_));
 XOR2x1_ASAP7_75t_R _1313_ (.A(net22),
    .Y(_0598_),
    .B(net8));
 NOR2x1_ASAP7_75t_R _1314_ (.A(net21),
    .B(_0421_),
    .Y(_0599_));
 AO221x1_ASAP7_75t_R _1315_ (.A1(net21),
    .A2(_0420_),
    .B1(_0598_),
    .B2(_0418_),
    .C(_0599_),
    .Y(_0731_));
 NAND2x1_ASAP7_75t_R _1316_ (.A(_0395_),
    .B(_0542_),
    .Y(_0600_));
 AND3x1_ASAP7_75t_R _1317_ (.A(_0404_),
    .B(_0395_),
    .C(_0542_),
    .Y(_0601_));
 AO21x1_ASAP7_75t_R _1318_ (.A1(_0391_),
    .A2(_0600_),
    .B(_0601_),
    .Y(_0733_));
 XOR2x1_ASAP7_75t_R _1319_ (.A(net32),
    .Y(_0602_),
    .B(net8));
 NOR2x1_ASAP7_75t_R _1320_ (.A(net31),
    .B(_0421_),
    .Y(_0603_));
 AO221x1_ASAP7_75t_R _1321_ (.A1(net31),
    .A2(_0420_),
    .B1(_0602_),
    .B2(_0418_),
    .C(_0603_),
    .Y(_0737_));
 XOR2x1_ASAP7_75t_R _1322_ (.A(net33),
    .Y(_0604_),
    .B(net8));
 NOR2x1_ASAP7_75t_R _1323_ (.A(net32),
    .B(_0421_),
    .Y(_0605_));
 AO221x1_ASAP7_75t_R _1324_ (.A1(net32),
    .A2(_0420_),
    .B1(_0604_),
    .B2(_0418_),
    .C(_0605_),
    .Y(_0739_));
 XOR2x1_ASAP7_75t_R _1325_ (.A(net31),
    .Y(_0606_),
    .B(net8));
 NOR2x1_ASAP7_75t_R _1326_ (.A(net30),
    .B(_0421_),
    .Y(_0607_));
 AO221x1_ASAP7_75t_R _1327_ (.A1(net30),
    .A2(_0420_),
    .B1(_0606_),
    .B2(_0418_),
    .C(_0607_),
    .Y(_0741_));
 XOR2x1_ASAP7_75t_R _1328_ (.A(net28),
    .Y(_0608_),
    .B(net8));
 NOR2x1_ASAP7_75t_R _1329_ (.A(net27),
    .B(_0421_),
    .Y(_0609_));
 AO221x1_ASAP7_75t_R _1330_ (.A1(net27),
    .A2(_0420_),
    .B1(_0608_),
    .B2(_0418_),
    .C(_0609_),
    .Y(_0745_));
 XOR2x1_ASAP7_75t_R _1331_ (.A(net29),
    .Y(_0610_),
    .B(net8));
 NOR2x1_ASAP7_75t_R _1332_ (.A(net28),
    .B(_0421_),
    .Y(_0611_));
 AO221x1_ASAP7_75t_R _1333_ (.A1(net28),
    .A2(_0420_),
    .B1(_0610_),
    .B2(_0418_),
    .C(_0611_),
    .Y(_0747_));
 XOR2x1_ASAP7_75t_R _1334_ (.A(net27),
    .Y(_0612_),
    .B(net8));
 NOR2x1_ASAP7_75t_R _1335_ (.A(net26),
    .B(_0421_),
    .Y(_0613_));
 AO221x1_ASAP7_75t_R _1336_ (.A1(net26),
    .A2(_0420_),
    .B1(_0612_),
    .B2(_0418_),
    .C(_0613_),
    .Y(_0749_));
 XOR2x1_ASAP7_75t_R _1337_ (.A(net26),
    .Y(_0614_),
    .B(net8));
 NOR2x1_ASAP7_75t_R _1338_ (.A(net25),
    .B(_0421_),
    .Y(_0615_));
 AO221x2_ASAP7_75t_R _1339_ (.A1(net25),
    .A2(_0420_),
    .B1(_0614_),
    .B2(_0418_),
    .C(_0615_),
    .Y(_0720_));
 XOR2x1_ASAP7_75t_R _1340_ (.A(net24),
    .Y(_0616_),
    .B(net8));
 NOR2x1_ASAP7_75t_R _1341_ (.A(net23),
    .B(_0421_),
    .Y(_0617_));
 AO221x1_ASAP7_75t_R _1342_ (.A1(net23),
    .A2(_0420_),
    .B1(_0616_),
    .B2(_0418_),
    .C(_0617_),
    .Y(_0751_));
 OA211x2_ASAP7_75t_R _1343_ (.A1(net169),
    .A2(net7),
    .B(_0372_),
    .C(net24),
    .Y(_0618_));
 INVx1_ASAP7_75t_R _1344_ (.A(_0618_),
    .Y(_0619_));
 OAI21x1_ASAP7_75t_R _1345_ (.A1(net24),
    .A2(_0705_),
    .B(_0619_),
    .Y(_0752_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 NOR2x2_ASAP7_75t_R _1347_ (.A(net1),
    .B(_0361_),
    .Y(_0621_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 OR3x1_ASAP7_75t_R _1349_ (.A(net84),
    .B(_0374_),
    .C(net174),
    .Y(_0623_));
 NOR2x1_ASAP7_75t_R _1350_ (.A(net171),
    .B(_0623_),
    .Y(_0624_));
 NOR2x2_ASAP7_75t_R _1351_ (.A(net1),
    .B(_0364_),
    .Y(_0625_));
 OA21x2_ASAP7_75t_R _1352_ (.A1(_0389_),
    .A2(_0623_),
    .B(_0625_),
    .Y(_0626_));
 AO21x1_ASAP7_75t_R _1353_ (.A1(_0621_),
    .A2(_0624_),
    .B(_0626_),
    .Y(_0084_));
 AND2x2_ASAP7_75t_R _1354_ (.A(_0414_),
    .B(net78),
    .Y(_0627_));
 NAND2x1_ASAP7_75t_R _1355_ (.A(net158),
    .B(_0627_),
    .Y(_0628_));
 AND3x1_ASAP7_75t_R _1356_ (.A(net158),
    .B(_0621_),
    .C(_0627_),
    .Y(_0629_));
 AO21x1_ASAP7_75t_R _1357_ (.A1(_0625_),
    .A2(_0628_),
    .B(_0629_),
    .Y(_0085_));
 AND3x2_ASAP7_75t_R _1358_ (.A(_0414_),
    .B(net78),
    .C(net174),
    .Y(_0630_));
 AND3x1_ASAP7_75t_R _1359_ (.A(_0411_),
    .B(_0621_),
    .C(_0630_),
    .Y(_0631_));
 AND4x1_ASAP7_75t_R _1360_ (.A(_0398_),
    .B(_0353_),
    .C(_0621_),
    .D(_0627_),
    .Y(_0632_));
 AND4x1_ASAP7_75t_R _1361_ (.A(net71),
    .B(_0398_),
    .C(_0405_),
    .D(_0627_),
    .Y(_0633_));
 OR2x4_ASAP7_75t_R _1362_ (.A(net1),
    .B(_0364_),
    .Y(_0634_));
 AOI211x1_ASAP7_75t_R _1363_ (.A1(_0411_),
    .A2(_0630_),
    .B(_0633_),
    .C(_0634_),
    .Y(_0635_));
 OR3x1_ASAP7_75t_R _1364_ (.A(_0631_),
    .B(_0632_),
    .C(_0635_),
    .Y(_0086_));
 INVx1_ASAP7_75t_R _1365_ (.A(_0627_),
    .Y(_0636_));
 NOR2x1_ASAP7_75t_R _1366_ (.A(_0401_),
    .B(_0636_),
    .Y(_0637_));
 OA21x2_ASAP7_75t_R _1367_ (.A1(_0401_),
    .A2(_0636_),
    .B(_0625_),
    .Y(_0638_));
 AO21x1_ASAP7_75t_R _1368_ (.A1(_0621_),
    .A2(_0637_),
    .B(_0638_),
    .Y(_0087_));
 OR3x1_ASAP7_75t_R _1369_ (.A(net84),
    .B(_0374_),
    .C(_0398_),
    .Y(_0639_));
 NOR2x1_ASAP7_75t_R _1370_ (.A(net171),
    .B(_0639_),
    .Y(_0640_));
 OA21x2_ASAP7_75t_R _1371_ (.A1(_0389_),
    .A2(_0639_),
    .B(_0625_),
    .Y(_0641_));
 AO21x1_ASAP7_75t_R _1372_ (.A1(_0621_),
    .A2(_0640_),
    .B(_0641_),
    .Y(_0088_));
 AND2x2_ASAP7_75t_R _1373_ (.A(net102),
    .B(net103),
    .Y(_0642_));
 AND2x4_ASAP7_75t_R _1374_ (.A(_0398_),
    .B(_0344_),
    .Y(_0643_));
 AO32x1_ASAP7_75t_R _1375_ (.A1(_0642_),
    .A2(_0537_),
    .A3(_0643_),
    .B1(_0630_),
    .B2(_0535_),
    .Y(_0644_));
 AOI221x1_ASAP7_75t_R _1376_ (.A1(_0535_),
    .A2(_0630_),
    .B1(_0643_),
    .B2(_0538_),
    .C(_0634_),
    .Y(_0645_));
 AO21x1_ASAP7_75t_R _1377_ (.A1(_0621_),
    .A2(_0644_),
    .B(_0645_),
    .Y(_0089_));
 AO32x1_ASAP7_75t_R _1378_ (.A1(net174),
    .A2(_0353_),
    .A3(_0627_),
    .B1(_0643_),
    .B2(_0411_),
    .Y(_0646_));
 AOI221x1_ASAP7_75t_R _1379_ (.A1(_0353_),
    .A2(_0630_),
    .B1(_0643_),
    .B2(_0411_),
    .C(_0634_),
    .Y(_0647_));
 AO21x1_ASAP7_75t_R _1380_ (.A1(_0621_),
    .A2(_0646_),
    .B(_0647_),
    .Y(_0090_));
 NAND2x1_ASAP7_75t_R _1381_ (.A(_0387_),
    .B(_0643_),
    .Y(_0648_));
 OR3x1_ASAP7_75t_R _1382_ (.A(net83),
    .B(_0642_),
    .C(_0426_),
    .Y(_0649_));
 OAI21x1_ASAP7_75t_R _1383_ (.A1(_0379_),
    .A2(_0648_),
    .B(_0649_),
    .Y(_0650_));
 OA211x2_ASAP7_75t_R _1384_ (.A1(_0379_),
    .A2(_0648_),
    .B(_0649_),
    .C(_0625_),
    .Y(_0651_));
 AO21x1_ASAP7_75t_R _1385_ (.A1(_0621_),
    .A2(_0650_),
    .B(_0651_),
    .Y(_0091_));
 NAND2x1_ASAP7_75t_R _1386_ (.A(_0398_),
    .B(_0344_),
    .Y(_0652_));
 NOR2x1_ASAP7_75t_R _1387_ (.A(net171),
    .B(_0652_),
    .Y(_0653_));
 OA21x2_ASAP7_75t_R _1388_ (.A1(_0389_),
    .A2(_0652_),
    .B(_0625_),
    .Y(_0654_));
 AO21x1_ASAP7_75t_R _1389_ (.A1(_0621_),
    .A2(_0653_),
    .B(_0654_),
    .Y(_0092_));
 NAND2x1_ASAP7_75t_R _1390_ (.A(_0344_),
    .B(net158),
    .Y(_0655_));
 AND3x1_ASAP7_75t_R _1391_ (.A(_0344_),
    .B(net158),
    .C(_0621_),
    .Y(_0656_));
 AO21x1_ASAP7_75t_R _1392_ (.A1(_0625_),
    .A2(_0655_),
    .B(_0656_),
    .Y(_0093_));
 AO32x1_ASAP7_75t_R _1393_ (.A1(net72),
    .A2(_0405_),
    .A3(_0643_),
    .B1(_0411_),
    .B2(_0345_),
    .Y(_0657_));
 AOI221x1_ASAP7_75t_R _1394_ (.A1(_0345_),
    .A2(_0411_),
    .B1(_0643_),
    .B2(_0353_),
    .C(_0634_),
    .Y(_0658_));
 AO21x1_ASAP7_75t_R _1395_ (.A1(_0621_),
    .A2(_0657_),
    .B(_0658_),
    .Y(_0094_));
 INVx1_ASAP7_75t_R _1396_ (.A(_0344_),
    .Y(_0659_));
 NOR2x1_ASAP7_75t_R _1397_ (.A(_0659_),
    .B(_0401_),
    .Y(_0660_));
 OA21x2_ASAP7_75t_R _1398_ (.A1(_0659_),
    .A2(_0401_),
    .B(_0625_),
    .Y(_0661_));
 AO21x1_ASAP7_75t_R _1399_ (.A1(_0621_),
    .A2(_0660_),
    .B(_0661_),
    .Y(_0095_));
 NAND2x1_ASAP7_75t_R _1400_ (.A(net174),
    .B(_0344_),
    .Y(_0662_));
 NOR2x1_ASAP7_75t_R _1401_ (.A(_0662_),
    .B(net171),
    .Y(_0663_));
 OA21x2_ASAP7_75t_R _1402_ (.A1(_0662_),
    .A2(net171),
    .B(_0625_),
    .Y(_0664_));
 AO21x1_ASAP7_75t_R _1403_ (.A1(_0621_),
    .A2(_0663_),
    .B(_0664_),
    .Y(_0096_));
 NAND2x1_ASAP7_75t_R _1404_ (.A(_0345_),
    .B(_0535_),
    .Y(_0665_));
 AND3x1_ASAP7_75t_R _1405_ (.A(_0345_),
    .B(_0535_),
    .C(_0621_),
    .Y(_0666_));
 AO21x1_ASAP7_75t_R _1406_ (.A1(_0625_),
    .A2(_0665_),
    .B(_0666_),
    .Y(_0097_));
 NOR2x1_ASAP7_75t_R _1407_ (.A(net1),
    .B(_0075_),
    .Y(_0098_));
 INVx5_ASAP7_75t_R _1408_ (.A(net1),
    .Y(_0667_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 AND2x2_ASAP7_75t_R _1410_ (.A(_0667_),
    .B(\add1.sm ),
    .Y(_0099_));
 AND2x2_ASAP7_75t_R _1411_ (.A(_0667_),
    .B(\ADDER.A1.Sum[0] ),
    .Y(_0100_));
 XOR2x1_ASAP7_75t_R _1412_ (.A(net89),
    .Y(_0669_),
    .B(_0038_));
 AND2x2_ASAP7_75t_R _1413_ (.A(_0667_),
    .B(_0669_),
    .Y(_0101_));
 OR3x1_ASAP7_75t_R _1414_ (.A(_0027_),
    .B(_0029_),
    .C(_0030_),
    .Y(_0670_));
 AND2x2_ASAP7_75t_R _1415_ (.A(_0449_),
    .B(_0670_),
    .Y(_0671_));
 XOR2x1_ASAP7_75t_R _1416_ (.A(net92),
    .Y(_0672_),
    .B(_0671_));
 AND2x2_ASAP7_75t_R _1417_ (.A(_0667_),
    .B(_0672_),
    .Y(_0102_));
 OA21x2_ASAP7_75t_R _1418_ (.A1(net91),
    .A2(_0671_),
    .B(_0039_),
    .Y(_0673_));
 XOR2x1_ASAP7_75t_R _1419_ (.A(net90),
    .Y(_0674_),
    .B(_0673_));
 AND2x2_ASAP7_75t_R _1420_ (.A(_0667_),
    .B(_0674_),
    .Y(_0103_));
 NOR2x1_ASAP7_75t_R _1421_ (.A(net1),
    .B(_0079_),
    .Y(_0104_));
 XNOR2x1_ASAP7_75t_R _1422_ (.B(_0078_),
    .Y(_0675_),
    .A(_0021_));
 AND2x2_ASAP7_75t_R _1423_ (.A(_0667_),
    .B(_0675_),
    .Y(_0105_));
 XOR2x1_ASAP7_75t_R _1424_ (.A(_0082_),
    .Y(_0676_),
    .B(_0454_));
 AND2x2_ASAP7_75t_R _1425_ (.A(_0667_),
    .B(_0676_),
    .Y(_0106_));
 OA21x2_ASAP7_75t_R _1426_ (.A1(_0082_),
    .A2(_0454_),
    .B(_0037_),
    .Y(_0677_));
 XOR2x1_ASAP7_75t_R _1427_ (.A(_0019_),
    .Y(_0678_),
    .B(_0677_));
 AND2x2_ASAP7_75t_R _1428_ (.A(_0667_),
    .B(_0678_),
    .Y(_0107_));
 NOR2x1_ASAP7_75t_R _1429_ (.A(net1),
    .B(_0077_),
    .Y(_0108_));
 XNOR2x1_ASAP7_75t_R _1430_ (.B(_0076_),
    .Y(_0679_),
    .A(_0015_));
 AND2x2_ASAP7_75t_R _1431_ (.A(_0667_),
    .B(_0679_),
    .Y(_0109_));
 XOR2x1_ASAP7_75t_R _1432_ (.A(_0012_),
    .Y(_0680_),
    .B(_0459_));
 AND2x2_ASAP7_75t_R _1433_ (.A(_0667_),
    .B(_0680_),
    .Y(_0110_));
 OA21x2_ASAP7_75t_R _1434_ (.A1(_0012_),
    .A2(_0459_),
    .B(_0036_),
    .Y(_0681_));
 XOR2x1_ASAP7_75t_R _1435_ (.A(_0013_),
    .Y(_0682_),
    .B(_0681_));
 AND2x2_ASAP7_75t_R _1436_ (.A(_0667_),
    .B(_0682_),
    .Y(_0111_));
 AND2x2_ASAP7_75t_R _1437_ (.A(\ADDER.A4.Sum[0] ),
    .B(_0667_),
    .Y(_0112_));
 XOR2x1_ASAP7_75t_R _1438_ (.A(_0032_),
    .Y(_0683_),
    .B(_0031_));
 AND2x2_ASAP7_75t_R _1439_ (.A(_0683_),
    .B(_0667_),
    .Y(_0113_));
 INVx2_ASAP7_75t_R _1440_ (.A(_0033_),
    .Y(_0684_));
 AO21x1_ASAP7_75t_R _1441_ (.A1(_0011_),
    .A2(_0460_),
    .B(_0010_),
    .Y(_0685_));
 AO21x1_ASAP7_75t_R _1442_ (.A1(_0081_),
    .A2(_0685_),
    .B(_0031_),
    .Y(_0686_));
 AND2x2_ASAP7_75t_R _1443_ (.A(_0034_),
    .B(_0686_),
    .Y(_0687_));
 XNOR2x1_ASAP7_75t_R _1444_ (.B(_0687_),
    .Y(_0688_),
    .A(_0684_));
 AND2x2_ASAP7_75t_R _1445_ (.A(_0667_),
    .B(_0688_),
    .Y(_0114_));
 AND3x1_ASAP7_75t_R _1446_ (.A(_0684_),
    .B(_0035_),
    .C(_0687_),
    .Y(_0689_));
 NOR2x1_ASAP7_75t_R _1447_ (.A(_0684_),
    .B(_0035_),
    .Y(_0690_));
 OA21x2_ASAP7_75t_R _1448_ (.A1(_0689_),
    .A2(_0690_),
    .B(_0667_),
    .Y(_0115_));
 INVx1_ASAP7_75t_R _1449_ (.A(_0030_),
    .Y(_0709_));
 INVx1_ASAP7_75t_R _1450_ (.A(_0727_),
    .Y(_0697_));
 FAx1_ASAP7_75t_R _1451_ (.SN(net101),
    .A(net166),
    .B(_0692_),
    .CI(_0693_),
    .CON(_0072_));
 FAx1_ASAP7_75t_R _1452_ (.SN(net88),
    .A(net100),
    .B(_0695_),
    .CI(_0696_),
    .CON(_0009_));
 FAx1_ASAP7_75t_R _1453_ (.SN(net163),
    .A(_0697_),
    .B(_0698_),
    .CI(_0699_),
    .CON(_0700_));
 FAx1_ASAP7_75t_R _1454_ (.SN(_0002_),
    .A(net87),
    .B(_0701_),
    .CI(_0702_),
    .CON(_0002_));
 FAx1_ASAP7_75t_R _1455_ (.SN(_0075_),
    .A(_0703_),
    .B(_0704_),
    .CI(_0705_),
    .CON(_0708_));
 FAx1_ASAP7_75t_R _1456_ (.SN(_0030_),
    .A(_0706_),
    .B(_0707_),
    .CI(_0708_),
    .CON(_0030_));
 FAx1_ASAP7_75t_R _1457_ (.SN(\ADDER.A4.Sum[0] ),
    .A(_0710_),
    .B(_0711_),
    .CI(_0712_),
    .CON(_0032_));
 FAx1_ASAP7_75t_R _1458_ (.SN(_0077_),
    .A(_0713_),
    .B(_0714_),
    .CI(_0715_),
    .CON(_0076_));
 FAx1_ASAP7_75t_R _1459_ (.SN(_0079_),
    .A(_0716_),
    .B(_0717_),
    .CI(_0451_),
    .CON(_0078_));
 FAx1_ASAP7_75t_R _1460_ (.SN(\ADDER.A1.Sum[0] ),
    .A(_0719_),
    .B(_0720_),
    .CI(_0709_),
    .CON(_0038_));
 HAxp5_ASAP7_75t_R _1461_ (.A(_0721_),
    .B(_0722_),
    .CON(_0727_),
    .SN(_0080_));
 HAxp5_ASAP7_75t_R _1462_ (.A(_0701_),
    .B(_0702_),
    .CON(_0000_),
    .SN(_0001_));
 HAxp5_ASAP7_75t_R _1463_ (.A(_0723_),
    .B(_0724_),
    .CON(_0005_),
    .SN(_0003_));
 HAxp5_ASAP7_75t_R _1464_ (.A(_0725_),
    .B(_0726_),
    .CON(_0006_),
    .SN(_0004_));
 HAxp5_ASAP7_75t_R _1465_ (.A(_0711_),
    .B(_0712_),
    .CON(_0081_),
    .SN(_0010_));
 HAxp5_ASAP7_75t_R _1466_ (.A(_0728_),
    .B(_0729_),
    .CON(_0036_),
    .SN(_0012_));
 HAxp5_ASAP7_75t_R _1467_ (.A(_0730_),
    .B(_0731_),
    .CON(_0011_),
    .SN(_0013_));
 HAxp5_ASAP7_75t_R _1468_ (.A(_0732_),
    .B(_0733_),
    .CON(_0014_),
    .SN(_0015_));
 HAxp5_ASAP7_75t_R _1469_ (.A(_0734_),
    .B(_0735_),
    .CON(_0016_),
    .SN(_0017_));
 HAxp5_ASAP7_75t_R _1470_ (.A(_0736_),
    .B(_0737_),
    .CON(_0037_),
    .SN(_0082_));
 HAxp5_ASAP7_75t_R _1471_ (.A(_0738_),
    .B(_0739_),
    .CON(_0018_),
    .SN(_0019_));
 HAxp5_ASAP7_75t_R _1472_ (.A(_0740_),
    .B(_0741_),
    .CON(_0020_),
    .SN(_0021_));
 HAxp5_ASAP7_75t_R _1473_ (.A(_0742_),
    .B(_0743_),
    .CON(_0022_),
    .SN(_0023_));
 HAxp5_ASAP7_75t_R _1474_ (.A(_0744_),
    .B(_0745_),
    .CON(_0039_),
    .SN(_0083_));
 HAxp5_ASAP7_75t_R _1475_ (.A(_0746_),
    .B(_0747_),
    .CON(_0024_),
    .SN(_0025_));
 HAxp5_ASAP7_75t_R _1476_ (.A(_0748_),
    .B(_0749_),
    .CON(_0026_),
    .SN(_0027_));
 HAxp5_ASAP7_75t_R _1477_ (.A(_0719_),
    .B(_0720_),
    .CON(_0028_),
    .SN(_0029_));
 HAxp5_ASAP7_75t_R _1478_ (.A(_0750_),
    .B(_0751_),
    .CON(_0034_),
    .SN(_0031_));
 HAxp5_ASAP7_75t_R _1479_ (.A(_0750_),
    .B(_0752_),
    .CON(_0035_),
    .SN(_0033_));
 DFFHQNx1_ASAP7_75t_R _1480_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0084_),
    .QN(_0071_));
 DFFHQNx3_ASAP7_75t_R _1481_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0085_),
    .QN(_0070_));
 DFFHQNx1_ASAP7_75t_R _1482_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0086_),
    .QN(_0069_));
 DFFHQNx3_ASAP7_75t_R _1483_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0087_),
    .QN(_0068_));
 DFFHQNx1_ASAP7_75t_R _1484_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0088_),
    .QN(_0067_));
 DFFHQNx1_ASAP7_75t_R _1485_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0089_),
    .QN(_0066_));
 DFFHQNx1_ASAP7_75t_R _1486_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0090_),
    .QN(_0065_));
 DFFHQNx3_ASAP7_75t_R _1487_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0091_),
    .QN(_0064_));
 DFFHQNx1_ASAP7_75t_R _1488_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0092_),
    .QN(_0063_));
 DFFHQNx3_ASAP7_75t_R _1489_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0093_),
    .QN(_0062_));
 DFFHQNx1_ASAP7_75t_R _1490_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0094_),
    .QN(_0061_));
 DFFHQNx1_ASAP7_75t_R _1491_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0095_),
    .QN(_0060_));
 DFFHQNx1_ASAP7_75t_R _1492_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0096_),
    .QN(_0059_));
 DFFHQNx3_ASAP7_75t_R _1493_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0097_),
    .QN(_0058_));
 DFFHQNx1_ASAP7_75t_R _1494_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0098_),
    .QN(_0057_));
 DFFHQNx1_ASAP7_75t_R _1495_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0099_),
    .QN(_0056_));
 DFFHQNx1_ASAP7_75t_R _1496_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0100_),
    .QN(_0055_));
 DFFHQNx1_ASAP7_75t_R _1497_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0101_),
    .QN(_0054_));
 DFFHQNx1_ASAP7_75t_R _1498_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0102_),
    .QN(_0053_));
 DFFHQNx1_ASAP7_75t_R _1499_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0103_),
    .QN(_0052_));
 DFFHQNx3_ASAP7_75t_R _1500_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0104_),
    .QN(_0051_));
 DFFHQNx1_ASAP7_75t_R _1501_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0105_),
    .QN(_0050_));
 DFFHQNx3_ASAP7_75t_R _1502_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0106_),
    .QN(_0049_));
 DFFHQNx1_ASAP7_75t_R _1503_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0107_),
    .QN(_0048_));
 DFFHQNx1_ASAP7_75t_R _1504_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0108_),
    .QN(_0047_));
 DFFHQNx3_ASAP7_75t_R _1505_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0109_),
    .QN(_0046_));
 DFFHQNx3_ASAP7_75t_R _1506_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0110_),
    .QN(_0045_));
 DFFHQNx3_ASAP7_75t_R _1507_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0111_),
    .QN(_0044_));
 DFFHQNx3_ASAP7_75t_R _1508_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0112_),
    .QN(_0043_));
 DFFHQNx3_ASAP7_75t_R _1509_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0113_),
    .QN(_0042_));
 DFFHQNx3_ASAP7_75t_R _1510_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0114_),
    .QN(_0041_));
 DFFHQNx3_ASAP7_75t_R _1511_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0115_),
    .QN(_0040_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Left_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Left_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Left_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Left_103 ();
 BUFx6f_ASAP7_75t_R input1 (.A(rst),
    .Y(net1));
 BUFx3_ASAP7_75t_R input2 (.A(x[0]),
    .Y(net2));
 BUFx6f_ASAP7_75t_R input3 (.A(x[10]),
    .Y(net3));
 BUFx6f_ASAP7_75t_R input4 (.A(x[11]),
    .Y(net4));
 BUFx12f_ASAP7_75t_R input5 (.A(x[12]),
    .Y(net5));
 BUFx6f_ASAP7_75t_R input6 (.A(x[13]),
    .Y(net6));
 BUFx4f_ASAP7_75t_R input7 (.A(x[14]),
    .Y(net7));
 BUFx16f_ASAP7_75t_R input8 (.A(x[15]),
    .Y(net8));
 BUFx3_ASAP7_75t_R input9 (.A(x[1]),
    .Y(net9));
 BUFx6f_ASAP7_75t_R input10 (.A(x[2]),
    .Y(net10));
 BUFx12f_ASAP7_75t_R input11 (.A(x[3]),
    .Y(net11));
 BUFx4f_ASAP7_75t_R input12 (.A(x[4]),
    .Y(net12));
 BUFx4f_ASAP7_75t_R input13 (.A(x[5]),
    .Y(net13));
 BUFx12f_ASAP7_75t_R input14 (.A(x[6]),
    .Y(net14));
 BUFx10_ASAP7_75t_R input15 (.A(x[7]),
    .Y(net15));
 BUFx3_ASAP7_75t_R input16 (.A(x[8]),
    .Y(net16));
 BUFx6f_ASAP7_75t_R input17 (.A(x[9]),
    .Y(net17));
 BUFx6f_ASAP7_75t_R input18 (.A(y[0]),
    .Y(net18));
 BUFx6f_ASAP7_75t_R input19 (.A(y[10]),
    .Y(net19));
 BUFx12_ASAP7_75t_R input20 (.A(y[11]),
    .Y(net20));
 BUFx6f_ASAP7_75t_R input21 (.A(y[12]),
    .Y(net21));
 BUFx4f_ASAP7_75t_R input22 (.A(y[13]),
    .Y(net22));
 BUFx10_ASAP7_75t_R input23 (.A(y[14]),
    .Y(net23));
 BUFx16f_ASAP7_75t_R input24 (.A(y[15]),
    .Y(net24));
 BUFx4f_ASAP7_75t_R input25 (.A(y[1]),
    .Y(net25));
 BUFx6f_ASAP7_75t_R input26 (.A(y[2]),
    .Y(net26));
 BUFx6f_ASAP7_75t_R input27 (.A(y[3]),
    .Y(net27));
 BUFx6f_ASAP7_75t_R input28 (.A(y[4]),
    .Y(net28));
 BUFx6f_ASAP7_75t_R input29 (.A(y[5]),
    .Y(net29));
 BUFx6f_ASAP7_75t_R input30 (.A(y[6]),
    .Y(net30));
 BUFx10_ASAP7_75t_R input31 (.A(y[7]),
    .Y(net31));
 BUFx4f_ASAP7_75t_R input32 (.A(y[8]),
    .Y(net32));
 BUFx6f_ASAP7_75t_R input33 (.A(y[9]),
    .Y(net33));
 BUFx2_ASAP7_75t_R output34 (.A(net34),
    .Y(p[0]));
 BUFx2_ASAP7_75t_R output35 (.A(net35),
    .Y(p[10]));
 BUFx2_ASAP7_75t_R output36 (.A(net36),
    .Y(p[11]));
 BUFx2_ASAP7_75t_R output37 (.A(net37),
    .Y(p[12]));
 BUFx2_ASAP7_75t_R output38 (.A(net38),
    .Y(p[13]));
 BUFx2_ASAP7_75t_R output39 (.A(net39),
    .Y(p[14]));
 BUFx2_ASAP7_75t_R output40 (.A(net40),
    .Y(p[15]));
 BUFx2_ASAP7_75t_R output41 (.A(net41),
    .Y(p[16]));
 BUFx2_ASAP7_75t_R output42 (.A(net42),
    .Y(p[17]));
 BUFx2_ASAP7_75t_R output43 (.A(net43),
    .Y(p[18]));
 BUFx2_ASAP7_75t_R output44 (.A(net44),
    .Y(p[19]));
 BUFx2_ASAP7_75t_R output45 (.A(net45),
    .Y(p[1]));
 BUFx2_ASAP7_75t_R output46 (.A(net46),
    .Y(p[20]));
 BUFx2_ASAP7_75t_R output47 (.A(net47),
    .Y(p[21]));
 BUFx2_ASAP7_75t_R output48 (.A(net48),
    .Y(p[22]));
 BUFx2_ASAP7_75t_R output49 (.A(net49),
    .Y(p[23]));
 BUFx2_ASAP7_75t_R output50 (.A(net50),
    .Y(p[24]));
 BUFx2_ASAP7_75t_R output51 (.A(net51),
    .Y(p[25]));
 BUFx2_ASAP7_75t_R output52 (.A(net52),
    .Y(p[26]));
 BUFx2_ASAP7_75t_R output53 (.A(net53),
    .Y(p[27]));
 BUFx2_ASAP7_75t_R output54 (.A(net54),
    .Y(p[28]));
 BUFx2_ASAP7_75t_R output55 (.A(net55),
    .Y(p[29]));
 BUFx2_ASAP7_75t_R output56 (.A(net56),
    .Y(p[2]));
 BUFx2_ASAP7_75t_R output57 (.A(net57),
    .Y(p[30]));
 BUFx2_ASAP7_75t_R output58 (.A(net58),
    .Y(p[31]));
 BUFx2_ASAP7_75t_R output59 (.A(net59),
    .Y(p[3]));
 BUFx2_ASAP7_75t_R output60 (.A(net60),
    .Y(p[4]));
 BUFx2_ASAP7_75t_R output61 (.A(net61),
    .Y(p[5]));
 BUFx2_ASAP7_75t_R output62 (.A(net62),
    .Y(p[6]));
 BUFx2_ASAP7_75t_R output63 (.A(net63),
    .Y(p[7]));
 BUFx2_ASAP7_75t_R output64 (.A(net64),
    .Y(p[8]));
 BUFx2_ASAP7_75t_R output65 (.A(net65),
    .Y(p[9]));
 BUFx4_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx4_ASAP7_75t_R clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_0__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_1__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_2__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_3__leaf_clk));
 BUFx2_ASAP7_75t_R rebuffer1 (.A(_0073_),
    .Y(net66));
 BUFx3_ASAP7_75t_R rebuffer2 (.A(net66),
    .Y(net67));
 BUFx2_ASAP7_75t_R rebuffer3 (.A(net67),
    .Y(net68));
 BUFx2_ASAP7_75t_R rebuffer4 (.A(net68),
    .Y(net69));
 BUFx2_ASAP7_75t_R rebuffer5 (.A(net68),
    .Y(net70));
 BUFx2_ASAP7_75t_R rebuffer6 (.A(net70),
    .Y(net71));
 BUFx2_ASAP7_75t_R rebuffer7 (.A(net71),
    .Y(net72));
 BUFx2_ASAP7_75t_R rebuffer8 (.A(net67),
    .Y(net73));
 BUFx2_ASAP7_75t_R rebuffer9 (.A(net73),
    .Y(net74));
 BUFx2_ASAP7_75t_R rebuffer10 (.A(net74),
    .Y(net75));
 BUFx2_ASAP7_75t_R rebuffer11 (.A(net73),
    .Y(net76));
 BUFx2_ASAP7_75t_R rebuffer12 (.A(_0074_),
    .Y(net77));
 BUFx2_ASAP7_75t_R rebuffer13 (.A(net77),
    .Y(net78));
 BUFx3_ASAP7_75t_R rebuffer14 (.A(net78),
    .Y(net79));
 BUFx2_ASAP7_75t_R rebuffer15 (.A(net79),
    .Y(net80));
 BUFx2_ASAP7_75t_R rebuffer16 (.A(net79),
    .Y(net81));
 BUFx6f_ASAP7_75t_R rebuffer17 (.A(net88),
    .Y(net82));
 BUFx2_ASAP7_75t_R rebuffer18 (.A(net82),
    .Y(net83));
 BUFx2_ASAP7_75t_R rebuffer19 (.A(net82),
    .Y(net84));
 BUFx2_ASAP7_75t_R rebuffer20 (.A(net88),
    .Y(net85));
 BUFx2_ASAP7_75t_R rebuffer21 (.A(net85),
    .Y(net86));
 BUFx2_ASAP7_75t_R rebuffer22 (.A(net164),
    .Y(net87));
 BUFx3_ASAP7_75t_R split23 (.A(_0009_),
    .Y(net88));
 BUFx2_ASAP7_75t_R rebuffer24 (.A(_0027_),
    .Y(net89));
 BUFx2_ASAP7_75t_R rebuffer25 (.A(_0025_),
    .Y(net90));
 BUFx2_ASAP7_75t_R rebuffer26 (.A(_0083_),
    .Y(net91));
 BUFx2_ASAP7_75t_R rebuffer27 (.A(net91),
    .Y(net92));
 BUFx4f_ASAP7_75t_R rebuffer28 (.A(_0389_),
    .Y(net93));
 BUFx2_ASAP7_75t_R rebuffer29 (.A(net93),
    .Y(net94));
 BUFx4f_ASAP7_75t_R rebuffer30 (.A(_0133_),
    .Y(net95));
 BUFx2_ASAP7_75t_R rebuffer31 (.A(net95),
    .Y(net96));
 BUFx2_ASAP7_75t_R rebuffer32 (.A(net95),
    .Y(net97));
 BUFx2_ASAP7_75t_R rebuffer33 (.A(net97),
    .Y(net98));
 BUFx2_ASAP7_75t_R rebuffer34 (.A(_0133_),
    .Y(net99));
 BUFx2_ASAP7_75t_R rebuffer35 (.A(net99),
    .Y(net100));
 BUFx2_ASAP7_75t_R split36 (.A(_0072_),
    .Y(net101));
 BUFx6f_ASAP7_75t_R rebuffer37 (.A(_0377_),
    .Y(net102));
 AO21x2_ASAP7_75t_R clone38 (.A1(_0346_),
    .A2(_0347_),
    .B(_0350_),
    .Y(net103));
 BUFx2_ASAP7_75t_R rebuffer90 (.A(_0170_),
    .Y(net155));
 BUFx2_ASAP7_75t_R rebuffer91 (.A(net155),
    .Y(net156));
 BUFx2_ASAP7_75t_R rebuffer92 (.A(net156),
    .Y(net157));
 BUFx2_ASAP7_75t_R rebuffer93 (.A(_0542_),
    .Y(net158));
 BUFx2_ASAP7_75t_R split94 (.A(net164),
    .Y(net159));
 BUFx2_ASAP7_75t_R split95 (.A(net164),
    .Y(net160));
 BUFx2_ASAP7_75t_R split96 (.A(net164),
    .Y(net161));
 BUFx2_ASAP7_75t_R split97 (.A(net164),
    .Y(net162));
 BUFx2_ASAP7_75t_R split98 (.A(net164),
    .Y(net163));
 BUFx3_ASAP7_75t_R rebuffer99 (.A(_0700_),
    .Y(net164));
 BUFx2_ASAP7_75t_R rebuffer100 (.A(_0171_),
    .Y(net165));
 BUFx2_ASAP7_75t_R rebuffer101 (.A(net165),
    .Y(net166));
 BUFx2_ASAP7_75t_R rebuffer102 (.A(_0183_),
    .Y(net167));
 BUFx2_ASAP7_75t_R rebuffer103 (.A(net167),
    .Y(net168));
 BUFx12_ASAP7_75t_R clone104 (.A(x[13]),
    .Y(net169));
 BUFx2_ASAP7_75t_R rebuffer105 (.A(_0131_),
    .Y(net170));
 OAI21x1_ASAP7_75t_R clone106 (.A1(_0379_),
    .A2(_0382_),
    .B(_0388_),
    .Y(net171));
 BUFx4f_ASAP7_75t_R clone107 (.A(x[13]),
    .Y(net172));
 BUFx2_ASAP7_75t_R rebuffer108 (.A(_0142_),
    .Y(net173));
 XNOR2x2_ASAP7_75t_R clone109 (.A(_0004_),
    .B(net101),
    .Y(net174));
 BUFx2_ASAP7_75t_R split110 (.A(_0002_),
    .Y(net175));
 BUFx8_ASAP7_75t_R clone111 (.A(x[13]),
    .Y(net176));
 BUFx2_ASAP7_75t_R rebuffer112 (.A(_0141_),
    .Y(net177));
 OR2x4_ASAP7_75t_R clone113 (.A(_0250_),
    .B(_0239_),
    .Y(net178));
 DECAPx10_ASAP7_75t_R FILLER_0_0_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_0_24 ();
 DECAPx2_ASAP7_75t_R FILLER_0_0_44 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_56 ();
 FILLER_ASAP7_75t_R FILLER_0_0_78 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_178 ();
 FILLER_ASAP7_75t_R FILLER_0_0_205 ();
 FILLER_ASAP7_75t_R FILLER_0_0_212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_219 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_241 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_24 ();
 FILLER_ASAP7_75t_R FILLER_0_1_36 ();
 FILLER_ASAP7_75t_R FILLER_0_1_44 ();
 FILLER_ASAP7_75t_R FILLER_0_1_52 ();
 FILLER_ASAP7_75t_R FILLER_0_1_64 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_76 ();
 FILLER_ASAP7_75t_R FILLER_0_1_87 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_92 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_158 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1_180 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_198 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_224 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1_246 ();
 FILLER_ASAP7_75t_R FILLER_0_1_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_262 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2 ();
 FILLER_ASAP7_75t_R FILLER_0_2_24 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_32 ();
 FILLER_ASAP7_75t_R FILLER_0_2_44 ();
 FILLER_ASAP7_75t_R FILLER_0_2_52 ();
 FILLER_ASAP7_75t_R FILLER_0_2_60 ();
 FILLER_ASAP7_75t_R FILLER_0_2_68 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_73 ();
 FILLER_ASAP7_75t_R FILLER_0_2_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_85 ();
 FILLER_ASAP7_75t_R FILLER_0_2_97 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_105 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_127 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_149 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_171 ();
 FILLER_ASAP7_75t_R FILLER_0_2_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_179 ();
 FILLER_ASAP7_75t_R FILLER_0_2_202 ();
 FILLER_ASAP7_75t_R FILLER_0_2_207 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_234 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_262 ();
 DECAPx4_ASAP7_75t_R FILLER_0_3_2 ();
 FILLER_ASAP7_75t_R FILLER_0_3_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_14 ();
 FILLER_ASAP7_75t_R FILLER_0_3_37 ();
 FILLER_ASAP7_75t_R FILLER_0_3_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_49 ();
 FILLER_ASAP7_75t_R FILLER_0_3_56 ();
 FILLER_ASAP7_75t_R FILLER_0_3_64 ();
 FILLER_ASAP7_75t_R FILLER_0_3_72 ();
 FILLER_ASAP7_75t_R FILLER_0_3_80 ();
 FILLER_ASAP7_75t_R FILLER_0_3_89 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_97 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_109 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_131 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_153 ();
 FILLER_ASAP7_75t_R FILLER_0_3_175 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_199 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_221 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_243 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_257 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_30 ();
 FILLER_ASAP7_75t_R FILLER_0_4_37 ();
 FILLER_ASAP7_75t_R FILLER_0_4_47 ();
 FILLER_ASAP7_75t_R FILLER_0_4_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_54 ();
 FILLER_ASAP7_75t_R FILLER_0_4_64 ();
 DECAPx1_ASAP7_75t_R FILLER_0_4_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_78 ();
 FILLER_ASAP7_75t_R FILLER_0_4_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_89 ();
 FILLER_ASAP7_75t_R FILLER_0_4_99 ();
 FILLER_ASAP7_75t_R FILLER_0_4_107 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_201 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_223 ();
 DECAPx6_ASAP7_75t_R FILLER_0_4_245 ();
 DECAPx1_ASAP7_75t_R FILLER_0_4_259 ();
 DECAPx2_ASAP7_75t_R FILLER_0_5_2 ();
 FILLER_ASAP7_75t_R FILLER_0_5_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_10 ();
 DECAPx6_ASAP7_75t_R FILLER_0_5_18 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_36 ();
 FILLER_ASAP7_75t_R FILLER_0_5_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_42 ();
 FILLER_ASAP7_75t_R FILLER_0_5_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_59 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_73 ();
 FILLER_ASAP7_75t_R FILLER_0_5_80 ();
 DECAPx2_ASAP7_75t_R FILLER_0_5_88 ();
 FILLER_ASAP7_75t_R FILLER_0_5_100 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_108 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_130 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_152 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_174 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_228 ();
 FILLER_ASAP7_75t_R FILLER_0_5_250 ();
 DECAPx2_ASAP7_75t_R FILLER_0_5_255 ();
 FILLER_ASAP7_75t_R FILLER_0_5_261 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_2 ();
 FILLER_ASAP7_75t_R FILLER_0_6_8 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_16 ();
 DECAPx4_ASAP7_75t_R FILLER_0_6_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_48 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_54 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_76 ();
 FILLER_ASAP7_75t_R FILLER_0_6_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_84 ();
 FILLER_ASAP7_75t_R FILLER_0_6_91 ();
 FILLER_ASAP7_75t_R FILLER_0_6_101 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_113 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_135 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_157 ();
 FILLER_ASAP7_75t_R FILLER_0_6_163 ();
 FILLER_ASAP7_75t_R FILLER_0_6_173 ();
 FILLER_ASAP7_75t_R FILLER_0_6_181 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_189 ();
 DECAPx4_ASAP7_75t_R FILLER_0_6_211 ();
 DECAPx4_ASAP7_75t_R FILLER_0_6_241 ();
 FILLER_ASAP7_75t_R FILLER_0_6_254 ();
 FILLER_ASAP7_75t_R FILLER_0_6_261 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_2 ();
 FILLER_ASAP7_75t_R FILLER_0_7_12 ();
 FILLER_ASAP7_75t_R FILLER_0_7_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_7_51 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_69 ();
 FILLER_ASAP7_75t_R FILLER_0_7_80 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_88 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_110 ();
 DECAPx2_ASAP7_75t_R FILLER_0_7_132 ();
 FILLER_ASAP7_75t_R FILLER_0_7_138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_7_150 ();
 FILLER_ASAP7_75t_R FILLER_0_7_156 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_164 ();
 FILLER_ASAP7_75t_R FILLER_0_7_176 ();
 DECAPx4_ASAP7_75t_R FILLER_0_7_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_194 ();
 FILLER_ASAP7_75t_R FILLER_0_7_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_203 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_210 ();
 DECAPx4_ASAP7_75t_R FILLER_0_7_234 ();
 FILLER_ASAP7_75t_R FILLER_0_7_247 ();
 FILLER_ASAP7_75t_R FILLER_0_7_254 ();
 FILLER_ASAP7_75t_R FILLER_0_7_261 ();
 FILLER_ASAP7_75t_R FILLER_0_8_2 ();
 FILLER_ASAP7_75t_R FILLER_0_8_11 ();
 DECAPx1_ASAP7_75t_R FILLER_0_8_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_26 ();
 FILLER_ASAP7_75t_R FILLER_0_8_35 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_43 ();
 DECAPx1_ASAP7_75t_R FILLER_0_8_55 ();
 DECAPx1_ASAP7_75t_R FILLER_0_8_71 ();
 DECAPx1_ASAP7_75t_R FILLER_0_8_83 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_96 ();
 DECAPx6_ASAP7_75t_R FILLER_0_8_118 ();
 FILLER_ASAP7_75t_R FILLER_0_8_132 ();
 FILLER_ASAP7_75t_R FILLER_0_8_141 ();
 DECAPx1_ASAP7_75t_R FILLER_0_8_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_162 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_169 ();
 FILLER_ASAP7_75t_R FILLER_0_8_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_177 ();
 DECAPx4_ASAP7_75t_R FILLER_0_8_184 ();
 FILLER_ASAP7_75t_R FILLER_0_8_194 ();
 FILLER_ASAP7_75t_R FILLER_0_8_204 ();
 DECAPx6_ASAP7_75t_R FILLER_0_8_212 ();
 FILLER_ASAP7_75t_R FILLER_0_8_226 ();
 FILLER_ASAP7_75t_R FILLER_0_8_234 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_262 ();
 DECAPx1_ASAP7_75t_R FILLER_0_9_2 ();
 FILLER_ASAP7_75t_R FILLER_0_9_14 ();
 FILLER_ASAP7_75t_R FILLER_0_9_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_26 ();
 FILLER_ASAP7_75t_R FILLER_0_9_47 ();
 FILLER_ASAP7_75t_R FILLER_0_9_55 ();
 DECAPx6_ASAP7_75t_R FILLER_0_9_61 ();
 FILLER_ASAP7_75t_R FILLER_0_9_75 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_83 ();
 FILLER_ASAP7_75t_R FILLER_0_9_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_91 ();
 DECAPx6_ASAP7_75t_R FILLER_0_9_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_111 ();
 DECAPx4_ASAP7_75t_R FILLER_0_9_119 ();
 FILLER_ASAP7_75t_R FILLER_0_9_134 ();
 FILLER_ASAP7_75t_R FILLER_0_9_152 ();
 FILLER_ASAP7_75t_R FILLER_0_9_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_168 ();
 DECAPx6_ASAP7_75t_R FILLER_0_9_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_191 ();
 FILLER_ASAP7_75t_R FILLER_0_9_206 ();
 FILLER_ASAP7_75t_R FILLER_0_9_215 ();
 FILLER_ASAP7_75t_R FILLER_0_9_223 ();
 DECAPx1_ASAP7_75t_R FILLER_0_9_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_235 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_262 ();
 FILLER_ASAP7_75t_R FILLER_0_10_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_4 ();
 FILLER_ASAP7_75t_R FILLER_0_10_11 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_27 ();
 DECAPx1_ASAP7_75t_R FILLER_0_10_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_39 ();
 DECAPx1_ASAP7_75t_R FILLER_0_10_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_62 ();
 FILLER_ASAP7_75t_R FILLER_0_10_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_70 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_83 ();
 FILLER_ASAP7_75t_R FILLER_0_10_89 ();
 FILLER_ASAP7_75t_R FILLER_0_10_96 ();
 DECAPx1_ASAP7_75t_R FILLER_0_10_103 ();
 DECAPx1_ASAP7_75t_R FILLER_0_10_127 ();
 FILLER_ASAP7_75t_R FILLER_0_10_138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_150 ();
 FILLER_ASAP7_75t_R FILLER_0_10_156 ();
 FILLER_ASAP7_75t_R FILLER_0_10_166 ();
 FILLER_ASAP7_75t_R FILLER_0_10_173 ();
 FILLER_ASAP7_75t_R FILLER_0_10_189 ();
 FILLER_ASAP7_75t_R FILLER_0_10_205 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_215 ();
 FILLER_ASAP7_75t_R FILLER_0_10_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_223 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_231 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_257 ();
 DECAPx4_ASAP7_75t_R FILLER_0_11_2 ();
 FILLER_ASAP7_75t_R FILLER_0_11_12 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_26 ();
 FILLER_ASAP7_75t_R FILLER_0_11_32 ();
 DECAPx1_ASAP7_75t_R FILLER_0_11_39 ();
 FILLER_ASAP7_75t_R FILLER_0_11_50 ();
 FILLER_ASAP7_75t_R FILLER_0_11_58 ();
 FILLER_ASAP7_75t_R FILLER_0_11_63 ();
 FILLER_ASAP7_75t_R FILLER_0_11_79 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_101 ();
 FILLER_ASAP7_75t_R FILLER_0_11_112 ();
 FILLER_ASAP7_75t_R FILLER_0_11_126 ();
 FILLER_ASAP7_75t_R FILLER_0_11_133 ();
 FILLER_ASAP7_75t_R FILLER_0_11_145 ();
 FILLER_ASAP7_75t_R FILLER_0_11_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_152 ();
 FILLER_ASAP7_75t_R FILLER_0_11_160 ();
 FILLER_ASAP7_75t_R FILLER_0_11_169 ();
 DECAPx4_ASAP7_75t_R FILLER_0_11_177 ();
 FILLER_ASAP7_75t_R FILLER_0_11_192 ();
 FILLER_ASAP7_75t_R FILLER_0_11_206 ();
 DECAPx1_ASAP7_75t_R FILLER_0_11_218 ();
 FILLER_ASAP7_75t_R FILLER_0_11_229 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_237 ();
 FILLER_ASAP7_75t_R FILLER_0_11_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_245 ();
 FILLER_ASAP7_75t_R FILLER_0_11_249 ();
 FILLER_ASAP7_75t_R FILLER_0_11_254 ();
 FILLER_ASAP7_75t_R FILLER_0_11_261 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_2 ();
 FILLER_ASAP7_75t_R FILLER_0_12_8 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_14 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_36 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_52 ();
 FILLER_ASAP7_75t_R FILLER_0_12_58 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_71 ();
 FILLER_ASAP7_75t_R FILLER_0_12_78 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_88 ();
 FILLER_ASAP7_75t_R FILLER_0_12_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_101 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_114 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_122 ();
 FILLER_ASAP7_75t_R FILLER_0_12_132 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_145 ();
 FILLER_ASAP7_75t_R FILLER_0_12_153 ();
 FILLER_ASAP7_75t_R FILLER_0_12_165 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_171 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_191 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_199 ();
 FILLER_ASAP7_75t_R FILLER_0_12_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_215 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_228 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_235 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_255 ();
 FILLER_ASAP7_75t_R FILLER_0_12_261 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_8 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_19 ();
 DECAPx4_ASAP7_75t_R FILLER_0_13_26 ();
 FILLER_ASAP7_75t_R FILLER_0_13_40 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_50 ();
 FILLER_ASAP7_75t_R FILLER_0_13_62 ();
 DECAPx4_ASAP7_75t_R FILLER_0_13_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_86 ();
 FILLER_ASAP7_75t_R FILLER_0_13_94 ();
 FILLER_ASAP7_75t_R FILLER_0_13_102 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_109 ();
 FILLER_ASAP7_75t_R FILLER_0_13_119 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_126 ();
 FILLER_ASAP7_75t_R FILLER_0_13_135 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_143 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_155 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_166 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_175 ();
 FILLER_ASAP7_75t_R FILLER_0_13_181 ();
 FILLER_ASAP7_75t_R FILLER_0_13_190 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_198 ();
 FILLER_ASAP7_75t_R FILLER_0_13_204 ();
 DECAPx4_ASAP7_75t_R FILLER_0_13_212 ();
 FILLER_ASAP7_75t_R FILLER_0_13_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_224 ();
 FILLER_ASAP7_75t_R FILLER_0_13_231 ();
 FILLER_ASAP7_75t_R FILLER_0_13_239 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_251 ();
 FILLER_ASAP7_75t_R FILLER_0_13_255 ();
 FILLER_ASAP7_75t_R FILLER_0_13_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_262 ();
 FILLER_ASAP7_75t_R FILLER_0_14_2 ();
 FILLER_ASAP7_75t_R FILLER_0_14_10 ();
 FILLER_ASAP7_75t_R FILLER_0_14_18 ();
 FILLER_ASAP7_75t_R FILLER_0_14_26 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_38 ();
 FILLER_ASAP7_75t_R FILLER_0_14_45 ();
 FILLER_ASAP7_75t_R FILLER_0_14_53 ();
 FILLER_ASAP7_75t_R FILLER_0_14_61 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_69 ();
 FILLER_ASAP7_75t_R FILLER_0_14_75 ();
 FILLER_ASAP7_75t_R FILLER_0_14_88 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_98 ();
 FILLER_ASAP7_75t_R FILLER_0_14_112 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_119 ();
 FILLER_ASAP7_75t_R FILLER_0_14_125 ();
 FILLER_ASAP7_75t_R FILLER_0_14_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_135 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_142 ();
 FILLER_ASAP7_75t_R FILLER_0_14_148 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_158 ();
 FILLER_ASAP7_75t_R FILLER_0_14_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_166 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_176 ();
 FILLER_ASAP7_75t_R FILLER_0_14_188 ();
 FILLER_ASAP7_75t_R FILLER_0_14_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_196 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_207 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_220 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_232 ();
 FILLER_ASAP7_75t_R FILLER_0_14_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_262 ();
 FILLER_ASAP7_75t_R FILLER_0_15_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_16 ();
 FILLER_ASAP7_75t_R FILLER_0_15_25 ();
 DECAPx2_ASAP7_75t_R FILLER_0_15_35 ();
 FILLER_ASAP7_75t_R FILLER_0_15_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_43 ();
 FILLER_ASAP7_75t_R FILLER_0_15_50 ();
 FILLER_ASAP7_75t_R FILLER_0_15_62 ();
 DECAPx6_ASAP7_75t_R FILLER_0_15_76 ();
 FILLER_ASAP7_75t_R FILLER_0_15_95 ();
 FILLER_ASAP7_75t_R FILLER_0_15_102 ();
 FILLER_ASAP7_75t_R FILLER_0_15_113 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_119 ();
 FILLER_ASAP7_75t_R FILLER_0_15_129 ();
 FILLER_ASAP7_75t_R FILLER_0_15_141 ();
 FILLER_ASAP7_75t_R FILLER_0_15_149 ();
 FILLER_ASAP7_75t_R FILLER_0_15_171 ();
 FILLER_ASAP7_75t_R FILLER_0_15_180 ();
 FILLER_ASAP7_75t_R FILLER_0_15_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_190 ();
 FILLER_ASAP7_75t_R FILLER_0_15_195 ();
 FILLER_ASAP7_75t_R FILLER_0_15_207 ();
 FILLER_ASAP7_75t_R FILLER_0_15_214 ();
 FILLER_ASAP7_75t_R FILLER_0_15_224 ();
 DECAPx2_ASAP7_75t_R FILLER_0_15_233 ();
 FILLER_ASAP7_75t_R FILLER_0_15_261 ();
 FILLER_ASAP7_75t_R FILLER_0_16_2 ();
 FILLER_ASAP7_75t_R FILLER_0_16_18 ();
 FILLER_ASAP7_75t_R FILLER_0_16_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_30 ();
 FILLER_ASAP7_75t_R FILLER_0_16_39 ();
 FILLER_ASAP7_75t_R FILLER_0_16_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_49 ();
 FILLER_ASAP7_75t_R FILLER_0_16_58 ();
 FILLER_ASAP7_75t_R FILLER_0_16_70 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_84 ();
 FILLER_ASAP7_75t_R FILLER_0_16_93 ();
 FILLER_ASAP7_75t_R FILLER_0_16_109 ();
 FILLER_ASAP7_75t_R FILLER_0_16_116 ();
 FILLER_ASAP7_75t_R FILLER_0_16_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_125 ();
 FILLER_ASAP7_75t_R FILLER_0_16_130 ();
 DECAPx1_ASAP7_75t_R FILLER_0_16_139 ();
 FILLER_ASAP7_75t_R FILLER_0_16_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_151 ();
 FILLER_ASAP7_75t_R FILLER_0_16_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_160 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_177 ();
 FILLER_ASAP7_75t_R FILLER_0_16_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_191 ();
 FILLER_ASAP7_75t_R FILLER_0_16_198 ();
 DECAPx1_ASAP7_75t_R FILLER_0_16_205 ();
 DECAPx1_ASAP7_75t_R FILLER_0_16_215 ();
 FILLER_ASAP7_75t_R FILLER_0_16_225 ();
 FILLER_ASAP7_75t_R FILLER_0_16_234 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_262 ();
 FILLER_ASAP7_75t_R FILLER_0_17_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_34 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_56 ();
 FILLER_ASAP7_75t_R FILLER_0_17_72 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_80 ();
 FILLER_ASAP7_75t_R FILLER_0_17_95 ();
 FILLER_ASAP7_75t_R FILLER_0_17_111 ();
 FILLER_ASAP7_75t_R FILLER_0_17_118 ();
 FILLER_ASAP7_75t_R FILLER_0_17_125 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_137 ();
 FILLER_ASAP7_75t_R FILLER_0_17_143 ();
 DECAPx4_ASAP7_75t_R FILLER_0_17_150 ();
 FILLER_ASAP7_75t_R FILLER_0_17_160 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_174 ();
 FILLER_ASAP7_75t_R FILLER_0_17_185 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_192 ();
 FILLER_ASAP7_75t_R FILLER_0_17_198 ();
 DECAPx6_ASAP7_75t_R FILLER_0_17_208 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_228 ();
 FILLER_ASAP7_75t_R FILLER_0_17_235 ();
 FILLER_ASAP7_75t_R FILLER_0_17_244 ();
 FILLER_ASAP7_75t_R FILLER_0_17_252 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_259 ();
 DECAPx2_ASAP7_75t_R FILLER_0_18_2 ();
 FILLER_ASAP7_75t_R FILLER_0_18_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_20 ();
 FILLER_ASAP7_75t_R FILLER_0_18_27 ();
 DECAPx4_ASAP7_75t_R FILLER_0_18_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_18_55 ();
 FILLER_ASAP7_75t_R FILLER_0_18_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_63 ();
 DECAPx6_ASAP7_75t_R FILLER_0_18_67 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_81 ();
 FILLER_ASAP7_75t_R FILLER_0_18_90 ();
 FILLER_ASAP7_75t_R FILLER_0_18_101 ();
 FILLER_ASAP7_75t_R FILLER_0_18_110 ();
 FILLER_ASAP7_75t_R FILLER_0_18_118 ();
 FILLER_ASAP7_75t_R FILLER_0_18_125 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_132 ();
 FILLER_ASAP7_75t_R FILLER_0_18_142 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_149 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_171 ();
 DECAPx6_ASAP7_75t_R FILLER_0_18_185 ();
 FILLER_ASAP7_75t_R FILLER_0_18_199 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_233 ();
 DECAPx2_ASAP7_75t_R FILLER_0_18_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_243 ();
 FILLER_ASAP7_75t_R FILLER_0_18_247 ();
 FILLER_ASAP7_75t_R FILLER_0_18_254 ();
 FILLER_ASAP7_75t_R FILLER_0_18_261 ();
 DECAPx2_ASAP7_75t_R FILLER_0_19_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_8 ();
 FILLER_ASAP7_75t_R FILLER_0_19_15 ();
 DECAPx4_ASAP7_75t_R FILLER_0_19_23 ();
 FILLER_ASAP7_75t_R FILLER_0_19_39 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_19_69 ();
 FILLER_ASAP7_75t_R FILLER_0_19_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_77 ();
 FILLER_ASAP7_75t_R FILLER_0_19_94 ();
 FILLER_ASAP7_75t_R FILLER_0_19_105 ();
 FILLER_ASAP7_75t_R FILLER_0_19_112 ();
 DECAPx4_ASAP7_75t_R FILLER_0_19_125 ();
 FILLER_ASAP7_75t_R FILLER_0_19_135 ();
 DECAPx2_ASAP7_75t_R FILLER_0_19_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_149 ();
 FILLER_ASAP7_75t_R FILLER_0_19_156 ();
 FILLER_ASAP7_75t_R FILLER_0_19_165 ();
 FILLER_ASAP7_75t_R FILLER_0_19_181 ();
 FILLER_ASAP7_75t_R FILLER_0_19_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_193 ();
 FILLER_ASAP7_75t_R FILLER_0_19_204 ();
 DECAPx2_ASAP7_75t_R FILLER_0_19_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_220 ();
 FILLER_ASAP7_75t_R FILLER_0_19_227 ();
 FILLER_ASAP7_75t_R FILLER_0_19_235 ();
 DECAPx2_ASAP7_75t_R FILLER_0_19_243 ();
 FILLER_ASAP7_75t_R FILLER_0_19_249 ();
 FILLER_ASAP7_75t_R FILLER_0_19_261 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_2 ();
 FILLER_ASAP7_75t_R FILLER_0_20_14 ();
 FILLER_ASAP7_75t_R FILLER_0_20_22 ();
 FILLER_ASAP7_75t_R FILLER_0_20_30 ();
 FILLER_ASAP7_75t_R FILLER_0_20_38 ();
 DECAPx6_ASAP7_75t_R FILLER_0_20_46 ();
 FILLER_ASAP7_75t_R FILLER_0_20_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_69 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_86 ();
 FILLER_ASAP7_75t_R FILLER_0_20_92 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_108 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_129 ();
 FILLER_ASAP7_75t_R FILLER_0_20_139 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_148 ();
 FILLER_ASAP7_75t_R FILLER_0_20_158 ();
 FILLER_ASAP7_75t_R FILLER_0_20_170 ();
 FILLER_ASAP7_75t_R FILLER_0_20_180 ();
 FILLER_ASAP7_75t_R FILLER_0_20_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_190 ();
 FILLER_ASAP7_75t_R FILLER_0_20_205 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_217 ();
 FILLER_ASAP7_75t_R FILLER_0_20_228 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_233 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_257 ();
 FILLER_ASAP7_75t_R FILLER_0_21_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_21_14 ();
 FILLER_ASAP7_75t_R FILLER_0_21_26 ();
 DECAPx1_ASAP7_75t_R FILLER_0_21_34 ();
 FILLER_ASAP7_75t_R FILLER_0_21_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_44 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_52 ();
 FILLER_ASAP7_75t_R FILLER_0_21_66 ();
 FILLER_ASAP7_75t_R FILLER_0_21_75 ();
 FILLER_ASAP7_75t_R FILLER_0_21_82 ();
 FILLER_ASAP7_75t_R FILLER_0_21_87 ();
 FILLER_ASAP7_75t_R FILLER_0_21_98 ();
 FILLER_ASAP7_75t_R FILLER_0_21_107 ();
 DECAPx6_ASAP7_75t_R FILLER_0_21_114 ();
 FILLER_ASAP7_75t_R FILLER_0_21_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_130 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_143 ();
 FILLER_ASAP7_75t_R FILLER_0_21_149 ();
 FILLER_ASAP7_75t_R FILLER_0_21_157 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_167 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_178 ();
 FILLER_ASAP7_75t_R FILLER_0_21_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_186 ();
 FILLER_ASAP7_75t_R FILLER_0_21_197 ();
 FILLER_ASAP7_75t_R FILLER_0_21_205 ();
 FILLER_ASAP7_75t_R FILLER_0_21_213 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_227 ();
 DECAPx1_ASAP7_75t_R FILLER_0_21_235 ();
 DECAPx1_ASAP7_75t_R FILLER_0_21_259 ();
 FILLER_ASAP7_75t_R FILLER_0_22_2 ();
 FILLER_ASAP7_75t_R FILLER_0_22_22 ();
 FILLER_ASAP7_75t_R FILLER_0_22_32 ();
 DECAPx1_ASAP7_75t_R FILLER_0_22_42 ();
 FILLER_ASAP7_75t_R FILLER_0_22_52 ();
 DECAPx4_ASAP7_75t_R FILLER_0_22_74 ();
 FILLER_ASAP7_75t_R FILLER_0_22_84 ();
 FILLER_ASAP7_75t_R FILLER_0_22_89 ();
 FILLER_ASAP7_75t_R FILLER_0_22_105 ();
 DECAPx1_ASAP7_75t_R FILLER_0_22_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_117 ();
 DECAPx4_ASAP7_75t_R FILLER_0_22_129 ();
 DECAPx4_ASAP7_75t_R FILLER_0_22_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_159 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_165 ();
 FILLER_ASAP7_75t_R FILLER_0_22_187 ();
 FILLER_ASAP7_75t_R FILLER_0_22_194 ();
 FILLER_ASAP7_75t_R FILLER_0_22_202 ();
 FILLER_ASAP7_75t_R FILLER_0_22_210 ();
 FILLER_ASAP7_75t_R FILLER_0_22_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_219 ();
 FILLER_ASAP7_75t_R FILLER_0_22_226 ();
 FILLER_ASAP7_75t_R FILLER_0_22_234 ();
 DECAPx1_ASAP7_75t_R FILLER_0_22_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_262 ();
 FILLER_ASAP7_75t_R FILLER_0_23_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_4 ();
 FILLER_ASAP7_75t_R FILLER_0_23_8 ();
 FILLER_ASAP7_75t_R FILLER_0_23_16 ();
 FILLER_ASAP7_75t_R FILLER_0_23_26 ();
 DECAPx4_ASAP7_75t_R FILLER_0_23_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_44 ();
 FILLER_ASAP7_75t_R FILLER_0_23_49 ();
 FILLER_ASAP7_75t_R FILLER_0_23_59 ();
 DECAPx6_ASAP7_75t_R FILLER_0_23_67 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_87 ();
 FILLER_ASAP7_75t_R FILLER_0_23_97 ();
 FILLER_ASAP7_75t_R FILLER_0_23_106 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_113 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_129 ();
 FILLER_ASAP7_75t_R FILLER_0_23_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_137 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_156 ();
 DECAPx6_ASAP7_75t_R FILLER_0_23_163 ();
 DECAPx4_ASAP7_75t_R FILLER_0_23_183 ();
 FILLER_ASAP7_75t_R FILLER_0_23_196 ();
 FILLER_ASAP7_75t_R FILLER_0_23_204 ();
 FILLER_ASAP7_75t_R FILLER_0_23_212 ();
 DECAPx4_ASAP7_75t_R FILLER_0_23_219 ();
 FILLER_ASAP7_75t_R FILLER_0_23_235 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_243 ();
 FILLER_ASAP7_75t_R FILLER_0_23_254 ();
 FILLER_ASAP7_75t_R FILLER_0_23_261 ();
 FILLER_ASAP7_75t_R FILLER_0_24_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_10 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_49 ();
 DECAPx4_ASAP7_75t_R FILLER_0_24_71 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_87 ();
 FILLER_ASAP7_75t_R FILLER_0_24_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_95 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_128 ();
 FILLER_ASAP7_75t_R FILLER_0_24_139 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_153 ();
 FILLER_ASAP7_75t_R FILLER_0_24_157 ();
 FILLER_ASAP7_75t_R FILLER_0_24_165 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_195 ();
 FILLER_ASAP7_75t_R FILLER_0_24_204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_212 ();
 DECAPx4_ASAP7_75t_R FILLER_0_24_234 ();
 FILLER_ASAP7_75t_R FILLER_0_24_244 ();
 FILLER_ASAP7_75t_R FILLER_0_24_249 ();
 FILLER_ASAP7_75t_R FILLER_0_24_254 ();
 FILLER_ASAP7_75t_R FILLER_0_24_261 ();
 FILLER_ASAP7_75t_R FILLER_0_25_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_10 ();
 DECAPx6_ASAP7_75t_R FILLER_0_25_32 ();
 FILLER_ASAP7_75t_R FILLER_0_25_46 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_51 ();
 FILLER_ASAP7_75t_R FILLER_0_25_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_59 ();
 DECAPx4_ASAP7_75t_R FILLER_0_25_68 ();
 FILLER_ASAP7_75t_R FILLER_0_25_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_80 ();
 DECAPx6_ASAP7_75t_R FILLER_0_25_91 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_109 ();
 DECAPx4_ASAP7_75t_R FILLER_0_25_116 ();
 FILLER_ASAP7_75t_R FILLER_0_25_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_128 ();
 DECAPx4_ASAP7_75t_R FILLER_0_25_138 ();
 FILLER_ASAP7_75t_R FILLER_0_25_148 ();
 FILLER_ASAP7_75t_R FILLER_0_25_156 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_166 ();
 FILLER_ASAP7_75t_R FILLER_0_25_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_174 ();
 FILLER_ASAP7_75t_R FILLER_0_25_181 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_189 ();
 FILLER_ASAP7_75t_R FILLER_0_25_195 ();
 FILLER_ASAP7_75t_R FILLER_0_25_204 ();
 FILLER_ASAP7_75t_R FILLER_0_25_212 ();
 DECAPx4_ASAP7_75t_R FILLER_0_25_220 ();
 FILLER_ASAP7_75t_R FILLER_0_25_230 ();
 FILLER_ASAP7_75t_R FILLER_0_25_252 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_257 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_26_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_38 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_46 ();
 FILLER_ASAP7_75t_R FILLER_0_26_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_68 ();
 DECAPx6_ASAP7_75t_R FILLER_0_26_90 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_110 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_121 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_128 ();
 FILLER_ASAP7_75t_R FILLER_0_26_134 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_150 ();
 FILLER_ASAP7_75t_R FILLER_0_26_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_158 ();
 FILLER_ASAP7_75t_R FILLER_0_26_165 ();
 FILLER_ASAP7_75t_R FILLER_0_26_173 ();
 FILLER_ASAP7_75t_R FILLER_0_26_181 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_189 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_201 ();
 FILLER_ASAP7_75t_R FILLER_0_26_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_209 ();
 DECAPx4_ASAP7_75t_R FILLER_0_26_217 ();
 FILLER_ASAP7_75t_R FILLER_0_26_233 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_245 ();
 FILLER_ASAP7_75t_R FILLER_0_26_249 ();
 FILLER_ASAP7_75t_R FILLER_0_26_254 ();
 FILLER_ASAP7_75t_R FILLER_0_26_261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_2 ();
 FILLER_ASAP7_75t_R FILLER_0_27_24 ();
 FILLER_ASAP7_75t_R FILLER_0_27_32 ();
 FILLER_ASAP7_75t_R FILLER_0_27_40 ();
 FILLER_ASAP7_75t_R FILLER_0_27_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_52 ();
 FILLER_ASAP7_75t_R FILLER_0_27_61 ();
 FILLER_ASAP7_75t_R FILLER_0_27_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_73 ();
 DECAPx1_ASAP7_75t_R FILLER_0_27_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_84 ();
 DECAPx4_ASAP7_75t_R FILLER_0_27_93 ();
 FILLER_ASAP7_75t_R FILLER_0_27_111 ();
 FILLER_ASAP7_75t_R FILLER_0_27_123 ();
 FILLER_ASAP7_75t_R FILLER_0_27_133 ();
 FILLER_ASAP7_75t_R FILLER_0_27_138 ();
 DECAPx4_ASAP7_75t_R FILLER_0_27_154 ();
 FILLER_ASAP7_75t_R FILLER_0_27_164 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_172 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_194 ();
 DECAPx1_ASAP7_75t_R FILLER_0_27_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_210 ();
 DECAPx1_ASAP7_75t_R FILLER_0_27_223 ();
 FILLER_ASAP7_75t_R FILLER_0_27_233 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_255 ();
 FILLER_ASAP7_75t_R FILLER_0_27_261 ();
 FILLER_ASAP7_75t_R FILLER_0_28_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_14 ();
 FILLER_ASAP7_75t_R FILLER_0_28_36 ();
 FILLER_ASAP7_75t_R FILLER_0_28_44 ();
 FILLER_ASAP7_75t_R FILLER_0_28_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_52 ();
 FILLER_ASAP7_75t_R FILLER_0_28_56 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_74 ();
 FILLER_ASAP7_75t_R FILLER_0_28_83 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_97 ();
 FILLER_ASAP7_75t_R FILLER_0_28_102 ();
 FILLER_ASAP7_75t_R FILLER_0_28_115 ();
 FILLER_ASAP7_75t_R FILLER_0_28_131 ();
 FILLER_ASAP7_75t_R FILLER_0_28_142 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_152 ();
 DECAPx6_ASAP7_75t_R FILLER_0_28_174 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_188 ();
 FILLER_ASAP7_75t_R FILLER_0_28_203 ();
 FILLER_ASAP7_75t_R FILLER_0_28_219 ();
 FILLER_ASAP7_75t_R FILLER_0_28_226 ();
 FILLER_ASAP7_75t_R FILLER_0_28_234 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_262 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_29_46 ();
 FILLER_ASAP7_75t_R FILLER_0_29_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_62 ();
 FILLER_ASAP7_75t_R FILLER_0_29_69 ();
 FILLER_ASAP7_75t_R FILLER_0_29_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_79 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_105 ();
 FILLER_ASAP7_75t_R FILLER_0_29_118 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_136 ();
 FILLER_ASAP7_75t_R FILLER_0_29_149 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_165 ();
 FILLER_ASAP7_75t_R FILLER_0_29_169 ();
 FILLER_ASAP7_75t_R FILLER_0_29_178 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_185 ();
 FILLER_ASAP7_75t_R FILLER_0_29_198 ();
 FILLER_ASAP7_75t_R FILLER_0_29_209 ();
 FILLER_ASAP7_75t_R FILLER_0_29_220 ();
 FILLER_ASAP7_75t_R FILLER_0_29_228 ();
 FILLER_ASAP7_75t_R FILLER_0_29_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_235 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_262 ();
 FILLER_ASAP7_75t_R FILLER_0_30_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_30_12 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_32 ();
 FILLER_ASAP7_75t_R FILLER_0_30_39 ();
 DECAPx1_ASAP7_75t_R FILLER_0_30_47 ();
 DECAPx4_ASAP7_75t_R FILLER_0_30_59 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_75 ();
 DECAPx6_ASAP7_75t_R FILLER_0_30_97 ();
 DECAPx1_ASAP7_75t_R FILLER_0_30_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_115 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_144 ();
 FILLER_ASAP7_75t_R FILLER_0_30_151 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_159 ();
 FILLER_ASAP7_75t_R FILLER_0_30_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_167 ();
 FILLER_ASAP7_75t_R FILLER_0_30_179 ();
 FILLER_ASAP7_75t_R FILLER_0_30_188 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_200 ();
 FILLER_ASAP7_75t_R FILLER_0_30_210 ();
 FILLER_ASAP7_75t_R FILLER_0_30_220 ();
 FILLER_ASAP7_75t_R FILLER_0_30_229 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_236 ();
 FILLER_ASAP7_75t_R FILLER_0_30_242 ();
 FILLER_ASAP7_75t_R FILLER_0_30_247 ();
 FILLER_ASAP7_75t_R FILLER_0_30_254 ();
 FILLER_ASAP7_75t_R FILLER_0_30_261 ();
 DECAPx6_ASAP7_75t_R FILLER_0_31_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_20 ();
 FILLER_ASAP7_75t_R FILLER_0_31_27 ();
 FILLER_ASAP7_75t_R FILLER_0_31_35 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_43 ();
 FILLER_ASAP7_75t_R FILLER_0_31_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_51 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_66 ();
 FILLER_ASAP7_75t_R FILLER_0_31_73 ();
 FILLER_ASAP7_75t_R FILLER_0_31_81 ();
 FILLER_ASAP7_75t_R FILLER_0_31_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_88 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_117 ();
 DECAPx6_ASAP7_75t_R FILLER_0_31_129 ();
 FILLER_ASAP7_75t_R FILLER_0_31_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_145 ();
 DECAPx4_ASAP7_75t_R FILLER_0_31_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_166 ();
 FILLER_ASAP7_75t_R FILLER_0_31_187 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_213 ();
 FILLER_ASAP7_75t_R FILLER_0_31_226 ();
 FILLER_ASAP7_75t_R FILLER_0_31_234 ();
 DECAPx4_ASAP7_75t_R FILLER_0_31_241 ();
 FILLER_ASAP7_75t_R FILLER_0_31_254 ();
 FILLER_ASAP7_75t_R FILLER_0_31_261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_24 ();
 FILLER_ASAP7_75t_R FILLER_0_32_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_32_40 ();
 FILLER_ASAP7_75t_R FILLER_0_32_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_66 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_79 ();
 FILLER_ASAP7_75t_R FILLER_0_32_87 ();
 FILLER_ASAP7_75t_R FILLER_0_32_97 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_105 ();
 FILLER_ASAP7_75t_R FILLER_0_32_121 ();
 DECAPx4_ASAP7_75t_R FILLER_0_32_129 ();
 FILLER_ASAP7_75t_R FILLER_0_32_151 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_163 ();
 FILLER_ASAP7_75t_R FILLER_0_32_174 ();
 DECAPx6_ASAP7_75t_R FILLER_0_32_182 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_202 ();
 FILLER_ASAP7_75t_R FILLER_0_32_211 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_229 ();
 FILLER_ASAP7_75t_R FILLER_0_32_236 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_262 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_24 ();
 FILLER_ASAP7_75t_R FILLER_0_33_36 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_51 ();
 DECAPx6_ASAP7_75t_R FILLER_0_33_62 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_80 ();
 FILLER_ASAP7_75t_R FILLER_0_33_87 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_101 ();
 DECAPx6_ASAP7_75t_R FILLER_0_33_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_137 ();
 FILLER_ASAP7_75t_R FILLER_0_33_150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_180 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_202 ();
 FILLER_ASAP7_75t_R FILLER_0_33_208 ();
 FILLER_ASAP7_75t_R FILLER_0_33_216 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_223 ();
 FILLER_ASAP7_75t_R FILLER_0_33_236 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_262 ();
 FILLER_ASAP7_75t_R FILLER_0_34_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_34_14 ();
 FILLER_ASAP7_75t_R FILLER_0_34_28 ();
 DECAPx1_ASAP7_75t_R FILLER_0_34_36 ();
 FILLER_ASAP7_75t_R FILLER_0_34_46 ();
 FILLER_ASAP7_75t_R FILLER_0_34_58 ();
 FILLER_ASAP7_75t_R FILLER_0_34_66 ();
 DECAPx1_ASAP7_75t_R FILLER_0_34_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_75 ();
 DECAPx4_ASAP7_75t_R FILLER_0_34_86 ();
 FILLER_ASAP7_75t_R FILLER_0_34_96 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_109 ();
 DECAPx6_ASAP7_75t_R FILLER_0_34_127 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_169 ();
 FILLER_ASAP7_75t_R FILLER_0_34_176 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_184 ();
 FILLER_ASAP7_75t_R FILLER_0_34_196 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_204 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_226 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_238 ();
 FILLER_ASAP7_75t_R FILLER_0_34_244 ();
 FILLER_ASAP7_75t_R FILLER_0_34_249 ();
 FILLER_ASAP7_75t_R FILLER_0_34_254 ();
 FILLER_ASAP7_75t_R FILLER_0_34_261 ();
 FILLER_ASAP7_75t_R FILLER_0_35_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_35_14 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_28 ();
 FILLER_ASAP7_75t_R FILLER_0_35_42 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_52 ();
 DECAPx4_ASAP7_75t_R FILLER_0_35_62 ();
 FILLER_ASAP7_75t_R FILLER_0_35_72 ();
 FILLER_ASAP7_75t_R FILLER_0_35_84 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_96 ();
 FILLER_ASAP7_75t_R FILLER_0_35_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_120 ();
 FILLER_ASAP7_75t_R FILLER_0_35_127 ();
 FILLER_ASAP7_75t_R FILLER_0_35_141 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_153 ();
 DECAPx4_ASAP7_75t_R FILLER_0_35_175 ();
 FILLER_ASAP7_75t_R FILLER_0_35_185 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_196 ();
 FILLER_ASAP7_75t_R FILLER_0_35_208 ();
 DECAPx6_ASAP7_75t_R FILLER_0_35_213 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_227 ();
 DECAPx6_ASAP7_75t_R FILLER_0_35_238 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_252 ();
 FILLER_ASAP7_75t_R FILLER_0_35_261 ();
 FILLER_ASAP7_75t_R FILLER_0_36_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_36_14 ();
 FILLER_ASAP7_75t_R FILLER_0_36_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_26 ();
 DECAPx4_ASAP7_75t_R FILLER_0_36_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_42 ();
 DECAPx6_ASAP7_75t_R FILLER_0_36_53 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_67 ();
 FILLER_ASAP7_75t_R FILLER_0_36_81 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_93 ();
 DECAPx4_ASAP7_75t_R FILLER_0_36_115 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_135 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_157 ();
 FILLER_ASAP7_75t_R FILLER_0_36_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_165 ();
 DECAPx6_ASAP7_75t_R FILLER_0_36_175 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_189 ();
 FILLER_ASAP7_75t_R FILLER_0_36_202 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_224 ();
 FILLER_ASAP7_75t_R FILLER_0_36_231 ();
 FILLER_ASAP7_75t_R FILLER_0_36_255 ();
 FILLER_ASAP7_75t_R FILLER_0_36_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_262 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_41 ();
 FILLER_ASAP7_75t_R FILLER_0_37_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_65 ();
 FILLER_ASAP7_75t_R FILLER_0_37_72 ();
 FILLER_ASAP7_75t_R FILLER_0_37_84 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_89 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_111 ();
 FILLER_ASAP7_75t_R FILLER_0_37_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_119 ();
 FILLER_ASAP7_75t_R FILLER_0_37_126 ();
 FILLER_ASAP7_75t_R FILLER_0_37_138 ();
 DECAPx6_ASAP7_75t_R FILLER_0_37_146 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_160 ();
 FILLER_ASAP7_75t_R FILLER_0_37_167 ();
 FILLER_ASAP7_75t_R FILLER_0_37_183 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_191 ();
 FILLER_ASAP7_75t_R FILLER_0_37_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_206 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_219 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_231 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_257 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_2 ();
 FILLER_ASAP7_75t_R FILLER_0_38_24 ();
 FILLER_ASAP7_75t_R FILLER_0_38_30 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_44 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_57 ();
 FILLER_ASAP7_75t_R FILLER_0_38_63 ();
 FILLER_ASAP7_75t_R FILLER_0_38_73 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_85 ();
 FILLER_ASAP7_75t_R FILLER_0_38_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_93 ();
 FILLER_ASAP7_75t_R FILLER_0_38_104 ();
 FILLER_ASAP7_75t_R FILLER_0_38_112 ();
 FILLER_ASAP7_75t_R FILLER_0_38_126 ();
 FILLER_ASAP7_75t_R FILLER_0_38_140 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_152 ();
 FILLER_ASAP7_75t_R FILLER_0_38_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_160 ();
 FILLER_ASAP7_75t_R FILLER_0_38_170 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_183 ();
 FILLER_ASAP7_75t_R FILLER_0_38_193 ();
 FILLER_ASAP7_75t_R FILLER_0_38_202 ();
 DECAPx6_ASAP7_75t_R FILLER_0_38_211 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_231 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_252 ();
 FILLER_ASAP7_75t_R FILLER_0_38_261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_2 ();
 FILLER_ASAP7_75t_R FILLER_0_39_24 ();
 DECAPx1_ASAP7_75t_R FILLER_0_39_38 ();
 FILLER_ASAP7_75t_R FILLER_0_39_52 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_69 ();
 FILLER_ASAP7_75t_R FILLER_0_39_78 ();
 DECAPx6_ASAP7_75t_R FILLER_0_39_88 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_112 ();
 FILLER_ASAP7_75t_R FILLER_0_39_134 ();
 FILLER_ASAP7_75t_R FILLER_0_39_142 ();
 DECAPx4_ASAP7_75t_R FILLER_0_39_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_164 ();
 FILLER_ASAP7_75t_R FILLER_0_39_171 ();
 FILLER_ASAP7_75t_R FILLER_0_39_185 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_194 ();
 DECAPx1_ASAP7_75t_R FILLER_0_39_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_216 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_224 ();
 FILLER_ASAP7_75t_R FILLER_0_39_230 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_238 ();
 FILLER_ASAP7_75t_R FILLER_0_39_244 ();
 FILLER_ASAP7_75t_R FILLER_0_39_249 ();
 FILLER_ASAP7_75t_R FILLER_0_39_254 ();
 FILLER_ASAP7_75t_R FILLER_0_39_261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_40_24 ();
 FILLER_ASAP7_75t_R FILLER_0_40_34 ();
 DECAPx1_ASAP7_75t_R FILLER_0_40_42 ();
 DECAPx6_ASAP7_75t_R FILLER_0_40_58 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_78 ();
 DECAPx4_ASAP7_75t_R FILLER_0_40_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_96 ();
 FILLER_ASAP7_75t_R FILLER_0_40_103 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_115 ();
 FILLER_ASAP7_75t_R FILLER_0_40_137 ();
 DECAPx4_ASAP7_75t_R FILLER_0_40_151 ();
 FILLER_ASAP7_75t_R FILLER_0_40_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_163 ();
 FILLER_ASAP7_75t_R FILLER_0_40_173 ();
 FILLER_ASAP7_75t_R FILLER_0_40_182 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_191 ();
 FILLER_ASAP7_75t_R FILLER_0_40_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_199 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_212 ();
 FILLER_ASAP7_75t_R FILLER_0_40_224 ();
 DECAPx1_ASAP7_75t_R FILLER_0_40_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_250 ();
 FILLER_ASAP7_75t_R FILLER_0_40_254 ();
 FILLER_ASAP7_75t_R FILLER_0_40_261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_24 ();
 FILLER_ASAP7_75t_R FILLER_0_41_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_32 ();
 FILLER_ASAP7_75t_R FILLER_0_41_39 ();
 DECAPx6_ASAP7_75t_R FILLER_0_41_51 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_71 ();
 FILLER_ASAP7_75t_R FILLER_0_41_80 ();
 FILLER_ASAP7_75t_R FILLER_0_41_90 ();
 FILLER_ASAP7_75t_R FILLER_0_41_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_100 ();
 FILLER_ASAP7_75t_R FILLER_0_41_113 ();
 DECAPx6_ASAP7_75t_R FILLER_0_41_121 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_139 ();
 FILLER_ASAP7_75t_R FILLER_0_41_146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_180 ();
 DECAPx6_ASAP7_75t_R FILLER_0_41_202 ();
 FILLER_ASAP7_75t_R FILLER_0_41_216 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_224 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_250 ();
 FILLER_ASAP7_75t_R FILLER_0_41_261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_42_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_37 ();
 DECAPx4_ASAP7_75t_R FILLER_0_42_59 ();
 FILLER_ASAP7_75t_R FILLER_0_42_69 ();
 FILLER_ASAP7_75t_R FILLER_0_42_79 ();
 FILLER_ASAP7_75t_R FILLER_0_42_84 ();
 FILLER_ASAP7_75t_R FILLER_0_42_98 ();
 FILLER_ASAP7_75t_R FILLER_0_42_107 ();
 FILLER_ASAP7_75t_R FILLER_0_42_119 ();
 DECAPx4_ASAP7_75t_R FILLER_0_42_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_137 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_150 ();
 FILLER_ASAP7_75t_R FILLER_0_42_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_174 ();
 FILLER_ASAP7_75t_R FILLER_0_42_184 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_193 ();
 FILLER_ASAP7_75t_R FILLER_0_42_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_201 ();
 DECAPx4_ASAP7_75t_R FILLER_0_42_208 ();
 FILLER_ASAP7_75t_R FILLER_0_42_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_226 ();
 FILLER_ASAP7_75t_R FILLER_0_42_249 ();
 FILLER_ASAP7_75t_R FILLER_0_42_254 ();
 FILLER_ASAP7_75t_R FILLER_0_42_261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_24 ();
 FILLER_ASAP7_75t_R FILLER_0_43_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_58 ();
 FILLER_ASAP7_75t_R FILLER_0_43_64 ();
 FILLER_ASAP7_75t_R FILLER_0_43_72 ();
 FILLER_ASAP7_75t_R FILLER_0_43_83 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_92 ();
 FILLER_ASAP7_75t_R FILLER_0_43_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_100 ();
 FILLER_ASAP7_75t_R FILLER_0_43_107 ();
 DECAPx6_ASAP7_75t_R FILLER_0_43_119 ();
 FILLER_ASAP7_75t_R FILLER_0_43_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_135 ();
 FILLER_ASAP7_75t_R FILLER_0_43_148 ();
 DECAPx6_ASAP7_75t_R FILLER_0_43_160 ();
 FILLER_ASAP7_75t_R FILLER_0_43_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_176 ();
 FILLER_ASAP7_75t_R FILLER_0_43_183 ();
 FILLER_ASAP7_75t_R FILLER_0_43_197 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_217 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_224 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_250 ();
 FILLER_ASAP7_75t_R FILLER_0_43_254 ();
 FILLER_ASAP7_75t_R FILLER_0_43_261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_30 ();
 FILLER_ASAP7_75t_R FILLER_0_44_35 ();
 FILLER_ASAP7_75t_R FILLER_0_44_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_44_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_65 ();
 FILLER_ASAP7_75t_R FILLER_0_44_72 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_80 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_116 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_144 ();
 DECAPx4_ASAP7_75t_R FILLER_0_44_151 ();
 FILLER_ASAP7_75t_R FILLER_0_44_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_163 ();
 FILLER_ASAP7_75t_R FILLER_0_44_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_175 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_182 ();
 FILLER_ASAP7_75t_R FILLER_0_44_204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_228 ();
 DECAPx4_ASAP7_75t_R FILLER_0_44_250 ();
 FILLER_ASAP7_75t_R FILLER_0_44_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_262 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_45_24 ();
 FILLER_ASAP7_75t_R FILLER_0_45_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_36 ();
 FILLER_ASAP7_75t_R FILLER_0_45_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_47 ();
 FILLER_ASAP7_75t_R FILLER_0_45_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_63 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_85 ();
 FILLER_ASAP7_75t_R FILLER_0_45_110 ();
 FILLER_ASAP7_75t_R FILLER_0_45_118 ();
 DECAPx4_ASAP7_75t_R FILLER_0_45_124 ();
 FILLER_ASAP7_75t_R FILLER_0_45_134 ();
 FILLER_ASAP7_75t_R FILLER_0_45_142 ();
 DECAPx6_ASAP7_75t_R FILLER_0_45_154 ();
 FILLER_ASAP7_75t_R FILLER_0_45_168 ();
 FILLER_ASAP7_75t_R FILLER_0_45_179 ();
 DECAPx2_ASAP7_75t_R FILLER_0_45_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_193 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_200 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_222 ();
 FILLER_ASAP7_75t_R FILLER_0_45_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_250 ();
 FILLER_ASAP7_75t_R FILLER_0_45_254 ();
 FILLER_ASAP7_75t_R FILLER_0_45_261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_46_24 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_38 ();
 DECAPx4_ASAP7_75t_R FILLER_0_46_50 ();
 FILLER_ASAP7_75t_R FILLER_0_46_60 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_65 ();
 FILLER_ASAP7_75t_R FILLER_0_46_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_73 ();
 DECAPx6_ASAP7_75t_R FILLER_0_46_84 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_98 ();
 FILLER_ASAP7_75t_R FILLER_0_46_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_112 ();
 FILLER_ASAP7_75t_R FILLER_0_46_120 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_128 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_146 ();
 FILLER_ASAP7_75t_R FILLER_0_46_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_154 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_163 ();
 FILLER_ASAP7_75t_R FILLER_0_46_173 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_195 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_227 ();
 DECAPx6_ASAP7_75t_R FILLER_0_46_249 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_47_24 ();
 FILLER_ASAP7_75t_R FILLER_0_47_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_36 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_43 ();
 FILLER_ASAP7_75t_R FILLER_0_47_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_59 ();
 FILLER_ASAP7_75t_R FILLER_0_47_69 ();
 FILLER_ASAP7_75t_R FILLER_0_47_77 ();
 FILLER_ASAP7_75t_R FILLER_0_47_87 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_95 ();
 FILLER_ASAP7_75t_R FILLER_0_47_105 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_121 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_133 ();
 FILLER_ASAP7_75t_R FILLER_0_47_140 ();
 FILLER_ASAP7_75t_R FILLER_0_47_153 ();
 FILLER_ASAP7_75t_R FILLER_0_47_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_163 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_173 ();
 FILLER_ASAP7_75t_R FILLER_0_47_189 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_197 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_225 ();
 DECAPx6_ASAP7_75t_R FILLER_0_47_247 ();
 FILLER_ASAP7_75t_R FILLER_0_47_261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_48_24 ();
 FILLER_ASAP7_75t_R FILLER_0_48_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_32 ();
 FILLER_ASAP7_75t_R FILLER_0_48_43 ();
 FILLER_ASAP7_75t_R FILLER_0_48_54 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_64 ();
 FILLER_ASAP7_75t_R FILLER_0_48_78 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_90 ();
 FILLER_ASAP7_75t_R FILLER_0_48_101 ();
 DECAPx4_ASAP7_75t_R FILLER_0_48_111 ();
 FILLER_ASAP7_75t_R FILLER_0_48_131 ();
 FILLER_ASAP7_75t_R FILLER_0_48_145 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_161 ();
 FILLER_ASAP7_75t_R FILLER_0_48_171 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_179 ();
 DECAPx2_ASAP7_75t_R FILLER_0_48_190 ();
 FILLER_ASAP7_75t_R FILLER_0_48_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_198 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_221 ();
 DECAPx6_ASAP7_75t_R FILLER_0_48_243 ();
 DECAPx2_ASAP7_75t_R FILLER_0_48_257 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_24 ();
 FILLER_ASAP7_75t_R FILLER_0_49_30 ();
 FILLER_ASAP7_75t_R FILLER_0_49_38 ();
 FILLER_ASAP7_75t_R FILLER_0_49_51 ();
 FILLER_ASAP7_75t_R FILLER_0_49_60 ();
 FILLER_ASAP7_75t_R FILLER_0_49_69 ();
 FILLER_ASAP7_75t_R FILLER_0_49_79 ();
 FILLER_ASAP7_75t_R FILLER_0_49_88 ();
 FILLER_ASAP7_75t_R FILLER_0_49_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_98 ();
 FILLER_ASAP7_75t_R FILLER_0_49_105 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_117 ();
 FILLER_ASAP7_75t_R FILLER_0_49_131 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_151 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_172 ();
 FILLER_ASAP7_75t_R FILLER_0_49_185 ();
 FILLER_ASAP7_75t_R FILLER_0_49_209 ();
 FILLER_ASAP7_75t_R FILLER_0_49_217 ();
 FILLER_ASAP7_75t_R FILLER_0_49_222 ();
 FILLER_ASAP7_75t_R FILLER_0_49_227 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_232 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_254 ();
 FILLER_ASAP7_75t_R FILLER_0_49_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_262 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_50_24 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_38 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_72 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_83 ();
 DECAPx6_ASAP7_75t_R FILLER_0_50_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_101 ();
 FILLER_ASAP7_75t_R FILLER_0_50_108 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_117 ();
 DECAPx4_ASAP7_75t_R FILLER_0_50_135 ();
 FILLER_ASAP7_75t_R FILLER_0_50_167 ();
 FILLER_ASAP7_75t_R FILLER_0_50_179 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_187 ();
 FILLER_ASAP7_75t_R FILLER_0_50_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_195 ();
 FILLER_ASAP7_75t_R FILLER_0_50_218 ();
 FILLER_ASAP7_75t_R FILLER_0_50_223 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_230 ();
 DECAPx4_ASAP7_75t_R FILLER_0_50_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_262 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_51_24 ();
 FILLER_ASAP7_75t_R FILLER_0_51_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_40 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_47 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_73 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_77 ();
 FILLER_ASAP7_75t_R FILLER_0_51_99 ();
 FILLER_ASAP7_75t_R FILLER_0_51_109 ();
 FILLER_ASAP7_75t_R FILLER_0_51_119 ();
 FILLER_ASAP7_75t_R FILLER_0_51_131 ();
 FILLER_ASAP7_75t_R FILLER_0_51_147 ();
 FILLER_ASAP7_75t_R FILLER_0_51_171 ();
 FILLER_ASAP7_75t_R FILLER_0_51_183 ();
 FILLER_ASAP7_75t_R FILLER_0_51_195 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_203 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_214 ();
 FILLER_ASAP7_75t_R FILLER_0_51_223 ();
 FILLER_ASAP7_75t_R FILLER_0_51_230 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_237 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_259 ();
endmodule
